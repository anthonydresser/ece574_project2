`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fqR67s8cBy/jbTeN196DpIBrWP6p4S7KSN05JgotCa3DCQok9PHpESJ+/YLHnMMyfVgYu3wMYulS
KP/HOuKOPw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o2f3dkiR8+1URrsaFkNAXM8HKCsrRh7Sklc6YYRJzdPn803OFcwNwVYhAiEMEOIJg1X2/T1BTFui
EQHVCIO1VCJStauI6Q8S2fTEfSbCGGuhlpfWUvhI0fluVmKgzRXGSxAPfzqyEe5IOj2rwzAzUH+w
I3b+vGSxoVxUbGLho4o=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ad3ngiL9tir1+ET0s4S3c+66wahwIoOVYNaNS7rfCSvbfk2aPsU2XB63og9D1Bg2SAX2HS1BQP3j
tM8/wIjLaDyunyJe0pY3Vy/MM/fpwDOYJVu9969hFmFD+MKjWmgclI/zBXndfn3HroxBNJ5YqbWw
T15thS0zDy/kMUmQm5Hhk2FofTiKZfDwJV8qMOs+IPoHxa32u/A5H/GAlLbYSj3iKXMDwdX1qvMx
Y/wH/Wca8f1dMVlyNgkzE7heSVl+umU4imcINE9Qacy9ksyf46mM/SkHQVg8M9UEek35LLEeFt+I
FDFYvl4xwj9zXwa6o3hy3BjN/8PdN/dXT3nHmg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
17s30izSWEvAAgQv6Vh1FDrqsfTI6ntDPxRKHcyQC5iftYo778GlTYz8H+ZoqnbRpo4Rx9iJh9p+
faDV0wcwXzKoFudL9jIBKm+gYqfFEvkVVJxOAlF/jWjG2nF/VmEXgcx03HwRaHCNUzX7tGZCK7Sm
cgQAO//GQtSMc3uUvyg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ru/nQZrQMQoFSUTnxErYixiyU4ARIhOaWewtUIoITFUVgG9z+gMss2pnsjU/kUZ9RWEI12+FXVka
+gRYtVpCxIPUEsXDftLv17WDI1tjcj5fWaceTamezhm6KUczosnGz9+NwbFG5z/2igcDAy6nQkqh
V58et0XyT53zqrn13mIfMOozEcd9PQwsZNuQCbg9wSERwoxnPdBLEg5UXNHZ0s6ahlbNehvtbbgl
yyf6RAnPelMgF4kT2YNl8xE5TPA5Ftff9vYHl3maAuj8YQ9wGLdONKEnZno1f+5yR5ljo2CbWnO+
oSovhdK1JX9QEbIkJ2QqxqDve6XKaLZUt7uHvQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NF2iKYemPHtuWn5hnoRCuPNs4c5eCM1mW9ddVILQydQ1OxFb70v0HA+tFCvBdEc/Oo23RE7HCPKv
BmrL9RcO1vKsdu91oZA6FdC/0KF7Iok4N8JN7IggHYwqedBTXbT1G79t+dcJQCYpp8IWyrFodnmv
7En+ptUiWn4gmkvJxLwkJl9miXUxtGBSTbY+MIpFl4u1hjtD6y8qRkjkITWWniMoIGON3+ShxVdH
vJ4+gC14V0VTb16Wd+kS1JZLUjkak6YQE2Y/wI+gM1SfXQv61yNCkzn4q8Fc5HhMXu8wvrAjPOoS
ZjZwz52Ph+N3YHEMsKW1FO0on8vy3THenmVVnQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`protect data_block
pa/mXep56TnCuXj5k+7cDUXVHoC8NVaoDetQOF7Qol+is+howENVqBnT9u3ujVh1MRLv7X/bo+Pw
dIaTRNqM13QI7LwDblH+oZidzWk5E+0o+q6XUe/PuIPWplhCAsUcdmA/8SXlHZ7izEXrMelk3K3E
hW31Yd8s2L8Q+jmE5ulzH5Ym2uefjH0z8D6P5t9Vv/wq3VtqEL9FzVpu8oNSX6URgx9B8xxnq01t
Fy0jYZrSGmZeJY9CWnoYYLHMO3+lU/rsKeQkM/S+ekNdfp7Iw98BhfwCgLE25GmXrWepjikkou9S
dKGZHUF+V21t18gZJQtRxiEGlzX4yjI6qhDlspAro92IvOSFv4YhatLnOiPU5/qzRyOv7lBh42f4
WnvEK92aaP4K3IKP9hUUQbZ6KbqtoA9Hu7Y6SHJaSgZdEcglsK41W40gL+4w9tcYftQDWGhazemk
Z2rjzkqfCStwishwyUC8HfuCd7vEomJrFQbZDp9UoEcwGW+KTunlUJdryCtTDByshGjMaG7pg63E
DU2pKgDNllOACA1p/M3P0RWfI0T1p9OUlkcdsYoGjwGHJINFPV75SDx2l1pN7UY/jOI0iuk8Gupk
7bGtBuhd4Xzdw6BoqqqQTxEl3msW1tHv296ggO7tRqP2MG6RDmZYnGQDWQ7bRaCjNDxOUZ3TInx0
weA1s0Ermeu0xznyXl/2cd5lXOxsAh8/NuRyp8gBhjVBQlM+XJ/ZN98pnMht+2A22ZV53PRRKWSI
md/nj5LSakYwBpVliQMJxKbpgj8ogI5941xc+TE7dnlHd6W95Z7s58RaXPcpSiOFwytY+2hdnJEJ
3kgLaoKonRQiyqsq7D04gwnqf4hgi+10N1Ceq7LqRYSokAPirdkgAPPqo9n8UGmq4A5Rq74ihl3o
lHoEr2IVZqlszpJNiFqkW0wv7OTrhER9KHLkaEIu7VVQAB4YY7EJjeyYgnF5Hgu1eOW91p9UgNph
Js+9XRLahOnFo+kAGB6RgrsZ2TTG853+qK+CUXBTT21+rU8gdLFdv496KOjTlluM4SiM4V/6o4uB
iETrxcNttSEF4Xeq1Cee1JTdUI62iR4a0NdV9NCjYtnFxDs1bxHZlk9oL+7ReHWzV7D8h87Dnpi6
0Rd9qRLJv+JOBufM66YiYbwlVjIkJ/R6HCdVcn99NrGb716K/1vF1x3t4VacZ2CbBZhiYJQf0K2M
kXkIjWejmpyux3/1FuGnTWsCwNeWBwftJIlKMpqa340lR5BM9OJPgnI28Hwq2YBQq3x+wKjLWhYz
1w8hjw11fIOoGppjkhOcDUIcTDQhKBiXxGgsE7Wupxc5NLAFqQ+WoBxjr+oN5TpZvN0MZO2mPmxG
rgPHNz8/+lYuG1FR8n9vSZUHJx8K48iVOAT/i14Y1o7xAa90xNAF8UFTK+H6ReWUWfNpbDiOHBKz
W8NmgrdJYtKj8lxHLNAPSrQaESojGl0Bt+Zq5N0CaxSyomg3Rf+jG+vYCPwPoFDS3TZroQ66Hr02
dJwzre7G1MYqQIqyPAjDbULPnE00AgM00b6XhOKFA9q4RIYVPqX4O2uJERi5LGHWCUzHxLUIZ/fT
SKpPJw7HC5mJ4IF1O2HaPmw1EHMI8T7JjOYkL1hN6LIuba50skH6GeEx+qJPVA3Dygyh8TduMDlh
YzP+XbomF5JLgDjEUTBbK3b8E1Z/JxFGUC3F4zyLUP+sL329FdP+eN+EdSJwlO5zQENsSsxfz7h5
Qi+Fdw3L95sUXAUlHpa3uavq/HCQ+u194RRdG9rFl5jrlE7/9eOjbaSdce665LJ+FvG3wKOFqbEd
Rn4DVNbll8NhvJgF0EA8FIbp5ARVQuu6tpMjPCMWz5wAAGaI7rY8B+b9WXglTeGd7EcrLZkIMnoK
0epw/9iwNKYD9ntlK6P6NFiLk8D7B9yuACAraUtXNwRFetpWz2us0uK8ROO6gHh+ab1wDNv8dMzM
TbImoCqc59vXKPbpyBNqCkQCBrbWRvfdPVkyOoeLkK6d/JBz5nbwq5zm/flsowu0MmTFplkA754W
TYgPckZ6Gw/OSy7Gl128KnOACPc+zuR+2I2XZePrTZoi/4mrM6aAtCzvRFw+JH6f2IeCPHgx2Uav
4dZDBv65z4rHF5UtrEfu5+tbXErnO1D4eVibaUJnud1fEVfxUDWSGkjejdZrASqNMU4E0Dc88aqf
fNbWty46dSk/0sGzJtz8j1ieTUErzBqUMj59fT52edQ9aWQuFeoubOCgOjAlahl6wNvs/6YrginB
92O9UlMA+Xr1h0XVtxcncF+Ivv1sz0lTg4gY3eke0G0xU8i1QYD1tfKnTQp9ltj0uBxIgFsWwJlm
8Mky65meLd0ZcnwB54xPLfca7I0MJ27OqEfyqCpYzupM5nCPzYn1bA+I4/njnkwWYK6gyNzgO0y6
zf4dfLMlfGT6lNggviTUpgZ45tEUQkAsKis//45qQB1y3rSbuBfeyQxYB2LYkmq+zUHR9g0grN+0
3Di5MoqpsvFgTbNgFQymjDqyT/FcQGAJu0jeDQ95RdnVLc2ksA7iEH6sIJPrWZMGqGZe8REpF8cX
ppz36viv8TplnNfHJZChB13fokYsMmYMDydN/8MI3XvxT0PD+WgEjamWd+pUikMZxk+ucRwrx+Ga
QvYTPbczD4cJP3yqWNSoRRqXcuS99+u8a4jgRvCTojLthBaI2iXL4eRyihtFHgzF102gKh8Zcyvp
V+TgZuvw3mBeteMnSrvvjfDKG9PTjW5c4mhZchjHb/mwOgooSLG229UeM1L4YmwRI+DFI7dw2r83
qin9aJ1xSwzd9qKWxpmCCBoo5Y2xfbUNIDk10VUqef9+NY2JGCiRcNcpE9LXquE0ooclN6flyDSM
V+vHaEur9BwUTisd9AINAtRlRKDCJ6Plt0Ld/1cZ0LZfKl4KTRqiuDGl+E5asfxLYUXBy6u0aRXw
WFo4jCQmg+ZwKrHrQ8H+dbsCTxqz0TndDpYbqqYmG0OUwBjOfd7v30dNCzqznkz681NhqGNG2Zgw
BcCLVFawpQ8cOaMPaJY5RXttak3kpZWx4EUzyiz0vRwkamsN0mT4hobQXVPFIUl9Gbhkqn8eu90p
yukhsKnCxEZE+VSsIj4DB3Y2zw1uo3GJPYx9RnAFws7Gn6aE3yW5SVUjNScvh1dCAijY299FQjPb
Y044uhHQJfJ4x/PlKgRi731/C320sWLTfKIlgPBERlWVaPG2ft4e4jCgtrkqeZLeEUpsF1NbwJBM
UdC1s5Uib1s3QbbqXhjnPEz1DZXQyJSSuQEQYsKfkI3RF4KxPPeAliIqLp8tYnUTeb+feWqA4LVC
C0Km37T10L1JVufz8BDh0/Gx1WzyD7vrq6IjKWRPL4XjDl9PMemDT7+OXzQ9wzdWAYJ1OboITCRP
405qcgbU+EaUsU+wwy04NWqg7Bdjd5gDjeDQDmzfDRF7drk+BsiA5JioiC8vU1xNKN2GmWMKPvvp
cf9nlNVg0BO8hd7sek8rgmdp+7sXjKzvMzEiFbSSbwNqRD9I74u2QpNM5Cr2nbeM40vLvt4RrCxP
lPNDIwS5JFFrlb6B4aBnE63RnlHHh+9WJ7WrIekMzyg1V0DkS5AvSH7zARTrmPGbUXEkG99AkWH0
dSIJCjlOwz1AUgGQRQz/lAX/KSgTDCVCssAcPKMXjxS1r8+jLjMmIklup13EOAyit0DWxHYSU4Vz
Svv+Xr3OCEjNxAOCtiWvk3+HgfR91oS/XnxeiQtG+nI+FNdXQ2LdW28za/y7kqkNE6vXz+q/RyD5
I5Y00nFb/bB+gd1+szn9EPMC9xdUwJqglEyZfQj9iremzJ3x202BxWWADf1J2RV2DFejtQtIuec6
4gPcgK+anuLx2D/41Oq8PasUJNcGltkkeIHCaRTjB6nhJ/Xcglhjq6JVJtUDfhv8LasbY01NMM68
F8a3aVEByQGbzOHSwrCeeUoWljeZMF2wefmwbtJeKW+wXx4pKYQMGTmyF5uFyXxYWf53Jx7gZGF3
ZFn9dLABjCZXYSBbtT9fzxgLLJFeEWvPfH/UM5kOj7rSLdNxGYUuZo0nbnvcSd+XokWggtL4auHs
Owme5Jbbiaf2gHWBprhE21Lvyyn7S4K7PyKjmR/d7N7e1TdMalQL/FetBYjG89hKZ4BfCkH13KGn
DRTDkM5+qDTl3ZPx4C8ZopGEyAv9zlSSPOQLUz8OwsF2lfOCczJVx7Y5vPqJP/SsaX9eLYvfxt+n
fm6DZ8Q8InqAETXG1Zv2/1Nk0WTkEjhimEBvyrfmzefRG5lYeOI7i2pvM9OAMIuaJh+Ct3vTusPO
DLSR3rAqrO+9eT6Nxjhi6gUcetrrAoGfiqEgiAv+mRWq2gsuO5Lv+xdpcjxqayEi9Av4OxAZXf9Q
gYqy0Svjo40CxRTbesGWovSbB8VMSBVrfvYme0Q3KGGT/eixbqRIxP2MlIH4hK8VTwSDneyZgopX
+jT54phXaGdLYu4kUsOf6akqpbQOdI2HoS8IWLP0LvZwrTfTwTRkftABYfKMvsteJlRclJ7kTdH+
gKE39KPubfY4psydKqd7ELSTGg/9mkIJIublLIXQzyoEcBw80RZOaLWGKajHNvbhZnBtov7JHlKD
pbq0tbIJgKaerZpAhauKnBEsuhROe75nWnet
`protect end_protected

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fqR67s8cBy/jbTeN196DpIBrWP6p4S7KSN05JgotCa3DCQok9PHpESJ+/YLHnMMyfVgYu3wMYulS
KP/HOuKOPw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o2f3dkiR8+1URrsaFkNAXM8HKCsrRh7Sklc6YYRJzdPn803OFcwNwVYhAiEMEOIJg1X2/T1BTFui
EQHVCIO1VCJStauI6Q8S2fTEfSbCGGuhlpfWUvhI0fluVmKgzRXGSxAPfzqyEe5IOj2rwzAzUH+w
I3b+vGSxoVxUbGLho4o=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ad3ngiL9tir1+ET0s4S3c+66wahwIoOVYNaNS7rfCSvbfk2aPsU2XB63og9D1Bg2SAX2HS1BQP3j
tM8/wIjLaDyunyJe0pY3Vy/MM/fpwDOYJVu9969hFmFD+MKjWmgclI/zBXndfn3HroxBNJ5YqbWw
T15thS0zDy/kMUmQm5Hhk2FofTiKZfDwJV8qMOs+IPoHxa32u/A5H/GAlLbYSj3iKXMDwdX1qvMx
Y/wH/Wca8f1dMVlyNgkzE7heSVl+umU4imcINE9Qacy9ksyf46mM/SkHQVg8M9UEek35LLEeFt+I
FDFYvl4xwj9zXwa6o3hy3BjN/8PdN/dXT3nHmg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
17s30izSWEvAAgQv6Vh1FDrqsfTI6ntDPxRKHcyQC5iftYo778GlTYz8H+ZoqnbRpo4Rx9iJh9p+
faDV0wcwXzKoFudL9jIBKm+gYqfFEvkVVJxOAlF/jWjG2nF/VmEXgcx03HwRaHCNUzX7tGZCK7Sm
cgQAO//GQtSMc3uUvyg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ru/nQZrQMQoFSUTnxErYixiyU4ARIhOaWewtUIoITFUVgG9z+gMss2pnsjU/kUZ9RWEI12+FXVka
+gRYtVpCxIPUEsXDftLv17WDI1tjcj5fWaceTamezhm6KUczosnGz9+NwbFG5z/2igcDAy6nQkqh
V58et0XyT53zqrn13mIfMOozEcd9PQwsZNuQCbg9wSERwoxnPdBLEg5UXNHZ0s6ahlbNehvtbbgl
yyf6RAnPelMgF4kT2YNl8xE5TPA5Ftff9vYHl3maAuj8YQ9wGLdONKEnZno1f+5yR5ljo2CbWnO+
oSovhdK1JX9QEbIkJ2QqxqDve6XKaLZUt7uHvQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NF2iKYemPHtuWn5hnoRCuPNs4c5eCM1mW9ddVILQydQ1OxFb70v0HA+tFCvBdEc/Oo23RE7HCPKv
BmrL9RcO1vKsdu91oZA6FdC/0KF7Iok4N8JN7IggHYwqedBTXbT1G79t+dcJQCYpp8IWyrFodnmv
7En+ptUiWn4gmkvJxLwkJl9miXUxtGBSTbY+MIpFl4u1hjtD6y8qRkjkITWWniMoIGON3+ShxVdH
vJ4+gC14V0VTb16Wd+kS1JZLUjkak6YQE2Y/wI+gM1SfXQv61yNCkzn4q8Fc5HhMXu8wvrAjPOoS
ZjZwz52Ph+N3YHEMsKW1FO0on8vy3THenmVVnQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 224608)
`protect data_block
pa/mXep56TnCuXj5k+7cDZsyudF/BgySsJRGxM0CTQyXaSNE43YiJ69HEvLxTJm8Ea4pTJ1v9WXi
nTRcVg9K3DHOhOIzICKejreObn6KOMYE3ly/M7H+fhzllYOKD5pk7B4yXp3+8guThANB+rWjHK9Y
QlXo/vrZRAqm5UugH2jL44bZl+J3MM6DOfPltMsaFdO80sD0MZ04Bl6G8KLijGLqxENyYwO0xYzX
NrELfVxNLtjvQbV+eijHqiV8Ce4D2pe88avTpBBsaA2LsNvF37qqgNO13VjqhnJ5ZKBsSYKaobTF
x2Ga70iOQOhT4OjBn9+U4pBJHZ4Wn5HPfMSX3sl85WeDA2h1ckeJ93XsxIrHtR7pzqDbcCQ95gR/
28mx16KCI5TXUkchCVx9ae9uYDsmuDY05eRcuZIHn5zR9GDnkk+Xn40C9ieTHKKramd/K74/P+Fg
u0vHnB+W3+xjbKeICuNWNxxBvq5gW/1Vl4USkW6pZhBF4SOyo7M17XxwnZyq4j1rbvNZLk9gIkPk
NNlwK6kE7B1L1H2uLuXIYHSVBT/OhLArS3yMoUxltu5XlLVY9PrXQjqVleqnUK4qpm6znhyExrJW
zFIrXUTh0og/6EEMDUGrr+zcEBCGvwl8DJs1p4SXxO1bbAP5RLJo0/8Xx++nzGSxszEutApZSVmc
uLv3O6QAmRMkNF7x71ZtX6beQOa0+4HbKd3+CMT0Wy8Q6szdQ7krEgJwsltJkPWbPbnB+n6yI5jq
Z0nQ+GrWJBZISyz9rq2Y42dHwivw19R3h2rJcOvCKRAhWSGYzVl/vYSzG2JxbN/OS02AbVNyUBhq
hIYJL801yH4KPTprDZbVdFFMvlXhr2MwRj0kay6mQwN5Yz7uBTQ/uGJYJumyW/fQqme67CZmu8Az
/593+kBJH1uy8fI9mTzneu9Z9Ab3+ylgooXP/QICiZATKXXjVofpko8qQlwkzbv0vNfolgbOfMO8
LGbPv/pko2E0drgqFc67Az9smYSdzLn9XGr0XVkK2To1R2GQ83mr3IyFyaaKqu9qlLGIOMP2L4Sy
VaxoXJ55/zKjbNp35rRNUC98eVbleNw3/bPxnVdFUP4cMcvFlRCGG5mqygeMLc6CoRvj7BGy9Zlf
+UlUDVvpzYRm/QbjUJ93LKBhF8h19pQSuUiLHXCac1YAvvpwY8yFF/ObDbkZ+q9ImDn/0DCV4i3r
Zrlmem7nqRKh9K/vnUM+KnUL13FTeyGc6LINYmOKX87BJNuPxXxaNYpEH0TvngWzpqtLnIj+NIAB
qgn3EZuAEsk0lHPzYZSeJWfbOCw04lumK7Xc7dCKWuTavFPFRrKtIne/8wyEV1t4PxJn1yj7y4Qc
LebsHACihr/ocajWb6ozhWKT6DNBsuCQmug+mi9xYaSxo/dlCWrgPWVEVQFBqPgHHJglqMGHJTcg
+UyQXBlGH/VJwqU2NewLdWfZPF09xqlOjARemreiabp8HDgx8gVTsjEsdYSrNjbBNSsyvDZ6bs75
YPrLUj8QX8j6+RPc9OMgaOupHpzhb8YW26bLGkqG0Ll8G++uaL/8GmhRD5OeW2OiWQapc6zRhhb9
0fwkX7LmFY46OrpZxpPznAhGbHmzjaDsn9B3dlhZ1pV9IIGrPyJS7v9lq64XzzXJ/pkbr6iTfKkK
HMu60seeskZGpgUK0BCdGoDi7ZRoee6aa2x/AyWBuUAhhx//jJQOSUlcXY0qLitL/dXV7KngWpJN
l4TJAPbguIi6GIqNVnBhOHPPvokMhKPWlIkZnOTbtNc/SweBkfyX7fA/+a7bmWb7d07puYv6nCsP
BQkNd7e9sExWb9EdXoy1MFBhWbN9PRVVlkt/k4z7MnKRn8NPQdoyYjg+19N2cO3qo3o6y41IR2oa
zjietIDYhP4KTANrala3HvdI92SNznP0X9Xu1PYizG5YiFSKrUS5FBXnbZtrUG7AuvNS5eA+P7Vk
5XGiTHXfdb2zvnAQ6Na2peNQDhCq7eZ2m+hGoRdd2eY8WBPd3lh18fJCPxYeqzfjznW+Dbe+oZXb
LTYAxMK5AF+Dy3exIcweB0UW7uiolShYeqFS2mrdYRVLWTdnWb1eUVwoCC6B353AVpWP0MHbizqA
iV1uglblL1pN7RitOGFVF367J1nCkWRW+cRrLUYnNik/7/7fhWIqbmiNxlP+tvx5SS5foO+uNATO
XVgnvVUOa1wrDNdBjcWTFg0VOMYUMs0bOHckn8LCmS+vvynSqbOmmwX+SnpKnBKavPyS6g5+H7Mw
C9iZy0E29GsOQCGagbLJsomYHyxf8SJTlmBEtS4oAcF+Fa44L50mrGGel/FkvfismVHtvqCflbL7
lJvttVdIR9UfV35Pt/M45fYayvbBulijzvpRWnmna7jFAUFb0KLIBZwWwcvIU2n8vY10SKI49X8/
LRJTuig/xDf/BkD3Ax5B6JzRwC2vwi/XxlfdlsviJvxfBcLduOy8r7bv4HlE1RaRmA16YBUqnmvV
27cLJT5tI9pzYP/zp6+E+EMIq2nxg9KVoJHLW+exjNLs2mGBw2c99Ji8YYDWOY2MQ7rpqzIItCBR
Tt8Rj03x8nL2v16qZbedESksXYsfz0yu5rKiHmGyv87DXVhPqgKr3sAWab3fcJR1DVCukKybu4h0
egy8AZpgwUV8TH8pgiU51bg1Al1AOb6K3parkkpttIfp8CVgHzZrxqcpPVyoe9hB/vBojp2tnTps
3yVGPxNmUfeSrRuk4XjpA1Ej2WxJGZ/zgDieHdWzHqUA8JLyfsJbMa/vpuClcFS5RwQnWna3mSZY
fW1J2Pq8SKYiqUt65Rnn/YUL4PCq9rG837qI2FsPozLe43mYaZwtgbh6B6yxfUALXmV+qUhsNQow
UC81q7R4bBUpo5d03gy+QNQEiyKqmaWSXI1ZYXCcfX1M0OR33KREDRj4HkgL6g+d84BgKKSiWcxP
/M1KDV1F+bjO+Xh4lRsIsbpAQA+QsTgVSX+4Uh5fZB9AatV9jACDw2wTpZrh0m4izQoV1KUaZpfL
LeGdhv/PQGtOIE6w/myalDA+KYWPujSDA8+Fit64kDlmVQGsb5xOm1NvUurix6d4uuK4APomKGlB
7SveS12xPybCZrI3HpxElVSOhWAHXlrNLHk8coU5ZVWAkyNwmLxp3vzquJYEttDmMsxtea58z8dF
+qKBLLguJ7H0g3FqOO5FCd2jip9jjeKCRMNw5EeRnxBWRurjcyT9ML06GEQLkewFG0QtAsM1+Oso
AuX+WapWsIEFiB+DvZAOjQBFnqvX2HAWX1kQT5aVMGqBUKQyp5VKYrz3kpKpIzQXuLCyfcIt+UpE
tEBTodYDQchY93ptRqxRKt7XResd3wRNsFzesF5tz2nXsEmhAEH219CKLPc81vcTyr4XqKk9UrFu
6PYmcWMUNIJ5ljsODBCjgYItb1Zdm4JevXG8w3MpeI7y2esDtG33H3nCBGajRnDBKoU697IM+FWR
4kODvCCzFy7q0xavnLStfpiASmFonMXhi7jbngzm72bwU4t+469Wo+pBOqNUp+P+H2jwafPSt6Ae
1flM2BHKpocj+9Iq0qPlAK481LvB2a1+IwuOMLu+kmZvEatWmXwU/dC7s8s43yWQPL/xh5Yjkt6k
gh7P2BBVevHLD5hNjjLF3N+3dZCS/wqxXVuioRTxqcAaKLdSv9hlDYQrd6aB4IhE/3spxO5JYfa6
x9bfGXuzzdL5YDO+2dha816seGE+OAUXogbBIop/f7yXGWI/9dvj8+MQjv6uU78azDk4r6MBhdzq
VhM2l70vYXdFnhkwcWhzRTIw+UgdAsjh/x8Rn56zqi4ql+/0zwZ5d3WD/Q3ZBWItwk/UQ2leQfjG
KZroUm9JzQd2uG7GaCXpX7Metr/oGufdQzYPlX1PJ/bTYueU635IB7Z1dRN4/RXuCjvcQmZIvgJ8
N7U3TIwZHypM3diLCzwvERbNdDlexZOwPhEZ4YHINUTIWuSKKuV3Y3DqBNUwFrrnA1gmaMoWEC+1
txXzDLnkThf0x36RYbVceTe9fh9oAWYKmo+EWuilODu4aUTnoYPei/tFMojDTQHShGNOVsVM02EG
NyJ/JjeqwodXcG+tZqVN2AZOfmQb1DQE5+GxvI5nDnpEmRVe6cU6HTsOwKt3r7dFWDSC7FZyi0CJ
x1aDKUZebQhOX3jYWv+Lxaq14MeWNI3bFxq8jViYzoy0R5sfbAPGQlOw/sTdM34X3aDW0AUNJzM0
zppk4EiRXG6ZdkvmJDxrfZx/h589h3jVYP1GkK5iLQ3czu0fnlWpI8l7bYP9sZ8CIdniHyxA5pUL
jxXZZJzS5AsIqS4gZaAgpY6jcLb/c9Hsl1E4jwqkA+vcmYSbue8LQYzmXJDnkg6PcBxPgdSf1MVk
i2BHZY+wHYSk4R+lRifYEO4iD3uwgK9Tnz6/rmW+Hoqnm0UnYu3bhhiog9pmpG4bbFlGR4zEVQ9G
DXQk34daXcW8LGljeZId6QqNTA2gMqpO9yLapLED41Jsua4CfIRPfiOfQ0uybTRq1oZM6l3gSj4n
2Y4NsciFEzuMObvpg2P8RWCfsDFGZgPPORKxLERLR/F2ob9oxnP4Ms0eAcvJqdBg60f/mbGe7NLB
T8yScsyjlutU//ayvcZwcKhgQ+hHJmWiBEDjB6++xScu+9RbC47PpYAR1Q2F6RC2WtUhcvqnkvPK
oBI5skXY79AmjAPtfUnEfs1v8MOO+BVvZVA6UDDIpAqy27nP5OgCT1fEL3ib/VwGLjo9a036LpLO
Yul/uQHS0+fN8wG1dOgPC4poNFQEPzz62z+Kj9rCHmoKtNvKnlFihqtKp+GULpV1H/Yy6TKdy/xn
NGAqVcj02yv/WihPzvpDurnw+WOLHWA/ItWmlxoCkNg8Zhau1S4U1Bvze0jcPyGalPtsMJt4zH/8
sLmi9dKcOlO8b76GWLD+XEzN9JvpoojeV0PTnBSbpjqNBcFkBMKEVxg1g3plZK6XQqycm7c4Qncv
lHpwe2ixgepiWyKxCnhfidhC3wT3T+ADmbXPBE84dZ9wyYVtWvz/tZCik/sHHpgoBrxyRmpnqJ6I
i8ePaCUZ6MPZcmwRtozc64XL0BAjY+R+vOGnJ/KSoj2tyW4AMKW8w55fgFdv9cDomJmi6ggZ8cus
xeikv1oPWdB1UTfSif9FYf/GVLIa5LNIGDpJ1UxeDNSMfcbNeD00DrTMdtAFh2QriLCwvJzKoIrB
oR1ZRVwbZnQMrMbAdAonpf3nIbJ0sIN3k/tI/KLr83DTkyprUrTfyrPOGOQfsbSYC6nVV4HUQBYH
KVcJIr0THUTAop/sdADDrApDngP8ipRyLBO+tw1t2Ux+BAJxpc7F/llLzMbKaiXJ7Yn0m2uIEFYn
i4LoPpdC/A4it6qcysT4SBTneGEB6y8No11VLju+YFXGbZJTeuHXcvw0EKrwTUYAUd5XAsua4zcb
T8s0QhYXKwKPgY0Hd00LlsAV/YCHKhn2x21NH0wqFfCbGGcbGSjzTEnaSOd6XCPc8p5zSLdZ9V+S
ob5nbtdTaNOEjpfE6kW6Xyb2lCRe/TpnpAFDJ6WGGn8MJOc9FzMitvHaWIm8tLApEmuMOyfbwE5q
K4y0vf8C5GnYtRTIG3DXQVCJwVFgMiyHh3yGYikTgJ3MuipogHdty3huGoFE6at8rRQiaCBaL/xf
zCUq6q5tH4oLlqEPviciYtKsmsLXCQ9t571jkKEto0Q1H+mI9HhhmWpm1Ts4I/k6HsO8zH2S23Q5
9UIGGoysBINPu5e0AFjN6mFsinBiEqTs2m3MwFpGHRnhosotjZsvtyzScaapJVrRG0dOgMtpEMZZ
V5611dFdub8Jqsix8563LkLIIAdVGhsB+q/jvMmUHhSmgM545jms1skbiBJu+hpN4AfxSWUaK3U/
b8QWWh/FBEDgV74K5TXWVyQn0uKH/327hoFWf3X26pu0V9nZx1k5aPXFQdPoEcmbXnxyEEUrei7r
DsJ4+IaahVUmj2vCr20noKg0e/fcriVh3hFTjtdWFGPpWMboHwsD71v3QjBwTB+UVMCQ5MwtnzGL
YFJU/bDIePm/Lq8cgDVAGWNrtBrEGDSfInXytwtJNfNo2yfmiKUFt3+O0OdmkBrt93mBn5IP2df1
HHS8JRjcCHgTb+n/62tfMPWTXmC5PRl5tFGqYn0vO+j/3uij+q66dOSFf7z4ow4VkSwmtSa0n6F1
xp5iPfhDx7lfdZnHtH4SWF6UJwrz/kPXtyLvulsPD1jSz6/lmZPOLldSKeTVdxj3WTOmjnqtAIm7
ltSAB9B7DIXOkCAeduD8muM3wYiFfEEKClVXSl5of+fx4pa488e10PgNRzKBIXH58z3Fysenrb0V
IVEXdcF118IdtJ2Y8n6D1rsubX93NzAMZfKqSlj7+h1c0mMqtgCUTJ4yXBYfPbo/xUzYGmPNeyRG
32pUaqgdZYt69+rS43FLhgK5pzPZldwr7RXcEv9gNY9Bqv8hCItiRq/GYnZyKky2g1TAwSh+y1ob
IaDZ4bd8RFriL88HX43qW8ReAsGMl6q+JlefcK4OjfUi9UKQHUtlov0D8yUDqff9iIQyFMpAs9uo
rPOQv4Bncyc5F+au3K/SmeoLHtFFXjIQIt86q8Erf6HLW7Ks9PUUnGZFJemLYiAByRD6+rhN/TlT
NaHn6j85jC0YYidlbb/kXpO237nORGhdJ0IfMsedUIFmRND+qM1oOYDrSFRSz+xzGGejmzdhip7l
dfDxXwDy5+UA/NKm1Y5tKAiK4KecjZr5cFpBSo4rCOJ4BPxg+ND3VRAA6GizDn7jFE8KOPvs5KcE
wvnObB49lZZHRDydnvTtDeQt2CNU67godbGvrWah2Q//P6MxgGxrwXywJQRGCOkthm6UQ74QGFjS
nUr0KEoeGeD+ZSF1oMdUkGbF9XAysUStOj1kjUn4fZPaVubcCkLtt6k53I4x76bsTyH9HPFahFxr
A2Qs/31jKaEMf09ohGHzrGCakeNCTHPTJvZpT+WoizSPQh5X0/Rsedf2f988qaynX5CLNCiar1GQ
DaSIW8HStdgPoLeAyKCY/32TRqFtjRstyC0TsT+d8p76+ig4P4CdCmGCDfJAWCzE44utMAdH3sIQ
tztkfhZ2aZ6x0ydy/mdtucF5hlB3K9u/cCkDZBVVrx6LBQA5EYFN9+jhXIMDq6CfVMhTy3L1c8M8
W+UETC3y2S0l9WO7KUKlpVKKFZLIz8RiWYYypJ/t8KV7f6K1ATOld9hcfM0Kj7mOEFRJ7wy9lmwF
J/BamGiCHGtjr6w13G028NPitk8iim5c/UUYbqTV2dEiL0fvtagkuqzt6zYtfkhdNEuARE/eZa/1
Cyib9WNjAjZFaPw6+yZpvFRBRv8ZxuOrO4KSPXT7fPVxZxLuE8Ay0O3M4vDSYkCei5a9vb0kiioJ
FQPVaNW+lUPmFgv+XyQHumluWDQE07iiNMeP0nzI9DJnMoAzjHGU9J/IY38b+fVLxY6KdXq7Mh+t
QrpkHtA9b47z/XGOaanZZ2gxXyGO21LzQd30K4jHHZqMD9QWxA6xL0Qx7zpGZb7muAFQbdXpPRmi
LCEH3Z2BW+roeDLYT4Zy99hXLK1OjQKoMoaLWBYx1Y+9tOLufcpCBitJ1+efN6urRjGctsOcIUkB
s2Dsy50WLWaEpSTj7473I1+NDUU2MbZy6sIZojGwXL6qtEVCtLh+uvyr57XClr/B+aGQ1nYsn51I
Yt/PSPKaOBWa7e7aqBFgeZAJRMWdsU0FfoSbTqJqUSAy4Z86VI0eBDBuroElxpcgy1bZV7WMvAtV
RjSQuYa0A7/L76j+rQ/yUd3JVLZB6Hh1H//T4JZu51B0SpRGXnICe9faCRjqatJXzV1ZFg4bZNcA
2OoEmoHub3w4dG/mcK55Lm7wLWbyqRsxhDiTtUeBoFLW0+YLsvEK7d/TXHCImcwIeslT/R/ZxY/q
VwcCSeHV3wsMPeTSRFoQsYrozx0u83gzF7qWzGA0dpQYO5LCFKwBzYCSiNpHSUfbSPdKp6YInNiJ
ncJqBMHq9Lm5h0wcMODg6NiXsARkNSSElIpQohW52kOyRz1C8RZaWKfL0WCKmvmFDqXqgPrbuNCa
fIaU4PzjJcqInSMkVKKemaT3LtUdo9FnemxnOWIcBen6UAnH3rLiMyahAsYQ1YypVY82CKqYMowQ
BZ/h80t8VoiEjxiMGMAAxMYVHEuZPbvRUnCq43a2GV93siMvVxnFWCd8vdCY2nIuXYT2jSycvhSd
zYzkLBxUOWmnhleddV4AiAOFHuk08mhuxWkuyWkmr+RfRfk/YMMTZEbAAI9xpepQUfFPcNdChLjk
KwWToTSMQQJNlmSi0pwOCIcqI+dUyPHWPaklfS4MSN5g79NT3/lhrZzQFo/xP+euKlc1GS/kROrJ
kBVkkvX4aV0zEiN82pP84hmYShSbGvutgwq7eEFEIfqfF24z+aAxCXlE463RzP92zAyEvPcgcnIt
Ihl7+L9GoY7r9HNoFixHUbmbxv3oIefEdxU6Jki8oXaBjARZfGJpNm3fOXe1jxEV5sFj3iamRVWg
8NBq/s8FdeIrG6JFGzhv8ECIgq56S8ygNsr87KCBHdNfVCn36D/WdJ3mymg+cQGvcdsCSnUIjIUd
656pz7PvHIuXYZ7o0K4FhCqEf9HitupPLBj4fPf582v4xM3TsyLC60i9L/NutgJYUWVfiNo9jURQ
LhR1Wpj9SOj6KQGhMD3pvPk/OzoQnL3uIZCJ6/imlUfVP07ylia82/cHAPQORMz7KIZCkonWxf3y
h6QiiauIWW74ZtJJHg4nuB+gm/J9PNUuhzpG6jaDTDsNoFo0RAEytnXMYkmU92zS95P91bbZCFZM
URN+fHPvZrHnd3nCk7Lr+4XZEZ/QHoDhu8e8IsBCD/6qB4Gs0RBzzttIjX3sgzKOsdvAMli9iktX
SuOZNbPDd9UCDnvLe3wdiYUhiDPeSqE/yNq+eNaZYB16/28D5MNRxBIxGcxGzSBX9mBR+6MdbMK7
j58+oWeJh/zxDfg3Edb0Q0VHajMYMchIrYLJB8ABHbajSz8rbvtashbKOArCXTYbu2I6e0UTwdNF
F7D4duqIpM1l3ilQtviUcoeTAfTWnVvkPm7ylnbt3jDOkXqGsRINiCQKeHjanN6uBPua8qma073P
8GeennMTPsdsOEB1F0L8IMC3gvUywb5nuYj5VoeLiSkZbibuuEATwNjNzwOgfHHX+e7nT+ajFdnn
CksZBjNqhYHyXEmbYAz1TnpC3Niqt4dHTO9cs0LTnThh70h02ugr/6a92G5PB9uKlfJtFFbPg2Dg
VXNcFks7uB+Y45QVTx5yjcNO0LnME7LwBfiipWe4aPCxA3dgfNi/rumRUELh71PTqdGJ1Mn9EhQn
owEXy9QGJ6ykKhwxhTlnZNrLP0bGNFCrw36K/f5yqshGSj36XcWLujRyv4xMXI2ql04ZFaKl8qfc
h/X1jiJZbAkxww80CQGh0lougxOUB7EHLcbKswftJ8X9dYfCvAKft7Yl8BJBeTqSQgQ2VlurGozW
VV4COV0aZgsVwMMxaoIKXoYZUzkOEX6Q2urMDdpdWe6+qU0FNlVdvwP0Uewrn3t6kf6bZ/b/SsTH
+Sy3y0CwLw1WaUdX+1sLpkPkv6rdMf41gnVqpAArANla2k8CzbSRGdlVezY1ln12PPw9Es4RTmnZ
JKXJXd2U4FCLiYwWs9KkxNyIFsdB4JTRvx8qQv4UrsK5Baf0XERYa+vZ1Cp5oqCI2R1DEjzw3r8k
OntrdxvpHX5HKLoBfTEfVo/dNZMVPKpmyBwBAYNcVd/VhB/11zo7TkniDdWKja6YT4qpSrBvM5bV
FfwCMT9sceFeoxRExOixD6cRZ+fNXfY+tBOep3ZvC9uo/+pqp7m6FyGNSN65ihgTqUbLPQZ8vvRd
O0RxU2tDP54RC/ZfDyWcKLq88hbDTVD1PByfV2YrQJCXH3YAXqRo67oul5B6dC6h9YrhV/7SpEcJ
kWg1IhWKg3/jBTPmDxs8UCiX2vsbSIoKSh1O6i5RltpV0SKHU3BNL67Pm1v0xnXzc13qo/QWw7cX
JL+Q/U65gT6zxfH3L6JLeWHcIzZEVStV2wkviXAcXVsxTPkEKaAkn4+fxecR4fjtz+t0lfCN2AxN
gxSs02JAb5AkfFVW2NCWNrwu+zqK7nSYVraKUTpOh89AiZyssthxcRBXY+N1idvf8ZGYa4wOtg7F
97ss+WdBhgqbI69F2to2mdxl9VdWjxVNuvN/6o2eAWAPI1W5iX60x0f7b+v591GSu8GraDqFdI8i
B0QlOyuLJdsYA2s7oodtDkR7uHth3hbB4p4ogv++z1gX9GrGmianX5fPTrekz+mzootG5ijMSmMA
AOSQIGfm4y3ZWrdENNC/IxEpDnahxspRoQnonmu5RPF9LcaMVIMqcOyPysLsuJMjWfEkaZ/HpIAe
wRgWwyN6Bornj5hEXBbuULE40O3SiC5JxEUoiaz/CLlUUPsEBxw+5m2xIxzcJbvA5IkBnLcSma5z
5E4cy62Y/PF1kNM0sQkXEqQPkrHt5HcCXGVWYHbTDur/T8ROVLEMQFg8LGrMvGbue8QpEod9c1gL
vEaMT9YKGY/BVLtTqCSf79bOvjiQ5IjK5CSRa4OawGLr2ywfYYTYsGLNWBMjRxH4Twmg2wStTx4B
1HObTm3zcxOycXPbqQUxNWUZryrSq1uhak7GD+fnenrxVFkD9Pv5h8+7qAb/fLuTR14+4w1rVkbX
vXaeE3rxRvd92iDqn/M8bNJeWkVD7lZ1TRVTzhaXy5yNRTlJ0n+2GJisyofzloGpRc0FYwC9GvXF
bzJoG8bmJiS3Zu1G8WrV3YnX/oxXWBQpvYqbtc5r8RdCgx0CNkX52RyKOYiCmm3I/6hCrzWguE53
L/CsFpVuhoSaNySnGDRMrJ3yUciM4ln8OQXw5wnu505Cikh+7hJhkBPwl2MJI7ma6Bf/+q4X92k5
1EJ4/IDp668UO1ufUQnzF8rlOH2LkjR9RWABFnIVs99xEB4oWmCtyYfmmVblOGwq3VxNE7QmPCcn
uwzzW06EZ5YdeJrgd48Cl3sC4WqG3tYuVNr5ZJVoY4o57gOUFinQUMQw3YWHIsc6I9SEuG/E4NFL
2TLWaXptmF3RxHCk5mY1EzVsRZCNBVUpdZkz4UlT1GQY5D5uDwIDo0l8tVKjCDUaK8XixSXYnx+T
n3k285wElp3RvOkqUh9tS4q3aQQpE5MkMNj+xpIrJ0HbQP2TOri5wM2REhzae7ElK8nlStUylLbJ
HU/H8hmRy1z35cSf2qOLska1JaBNaDv8s4C0C7ZOkqWGlNcGJWhqAe7RAM8VCOxI8vrpvebA7DGx
B9q/LaHvXlq5ViAq78I1NEqYDkBYDB3jXnzWhWQU03Gzj3CtTiYeXirhrTI9mGb93eyFR+1MUSv1
/wbKJQC6XXix52fxCPbMxh0OWutYBbb4+njvWNLTwZao3HNG141QH+J27vIgzw1B/GNVOZTTcW6x
9xJZFThWoVhNi/1avjSSlBuocalkTHXu7iO0B+k3cfA+QjoWgYPeMl8iOcga6Zpqx4CmvsMI2GdK
WaLV2YrhIMiGyQp0OM6IFWfE6tJ/Wtn6CzdDKvHGWm7dlZs0lVZXvS0il4rrSkB7I4iQt0Z9VZL5
rIU0AI3+5U4s8claYbXRap+MT2TPqxckPiTmFYOrPy04qCqfJjRdTe40RrIcVbb5EfuwETpBT/M4
YH4Jc/zRTqNtEGARV5/mx9WkrlD/P38eVO08wwSXtF+CRNiNFhGtcXUc43JppSFVL3vvMk8ZBbI5
zXrKTHZyDA8rXdtZOotaf8fRdDioVBdFTpwbsQ0c4Lybveq8dpA0kBSH3ytR6zJqzJycFw6y6D0R
yDIvBS0aQ93MPlRNu5dp1bT9Hs/18BiVPGR7Iel8XTYNnlusPwzuvnZ4BRs9VGUtNTtB3GTx7s/U
Dekg1ggyhSOWsn4d9WVOrAgvZ1MeWYlXsZkC8UFAH4apY9Dvj/OBcsgQhQ25IBpUIV7ZBknBmxRD
W5C8+WHo9rn9LVByed5ZZlsjzLKbRBaMiVbMH8HzFcOrhw7HJ9rEPluQz4LE7K/2dyzfDuZbD3uB
9NDl+7SlpMgk5PMNMC6ePGkgxcI5p24tfAbRE+3xRwxkW2cKJ1OOHZsfWAJXrAwDU8856yebFhAQ
qfQagodlhYb4C3phF5QGi5sZ/LcUMALQK7jDU7W2dPzOsZAmKqimU08ESJEyAM3aq0Zzj3K3Ade+
cOweNJos5dDvxDwxGrbI2cD/WaoE9mNo8mHI7NslPRZE32/OOwTpYarULgcrqm2npjWLv+RkyC4m
QNy7/BjinvYNrbwBL9l7GJOTzzYQqeVUqeEN9bLaY1Cw+nbtacj6cW+IwnFY7ELXWCgcrnTucnk1
e3iBn+JSMi9PK1d+V5kO2p5JQC/n5BxjNt2QZWv1syXAoC8Izs8vnf5aLqoNesV8lvfeZf1iJR0P
5PKDQVvfu03kpWovrXVPSo7zOdA7kMqGm7Hy68bgX0cV5XjFrgyeUJB2HbKgNqAHfhUSctAHEzyz
9NYZQvaeW7qNXy+/U13DyrlGBw5G+UzNC4kDyogRSH8oBOdcvRK802VyAGZQ0kf26eTf8AZnwrpl
LgYkp55KmUSkDlj+FaXeYD+yvJFLb8MpHHAJ/BZtq6jEbaOLc6WazuhdGeKFS5qyByiI2bxm5EZw
t098aE9R5YxCk2vJZnvrgVYj3nFZxZQAsl9pTtRNtT6KMLQFUhKVXvrl+QaY4jzmCJuegrFwYG0W
NvyJ9UCnf828657UGuF5FIqq5FS1ZPjlXvxK9QYD0KpdAMba2CHbwpmKocJZIdQQJiGVxJUao4ar
537mqN095LExxAo4fBE57ar2W0oOgiNY/0CvCDQVq9TVE//ErPLbju3yga9GtAa08T6yg491iAGu
Hx51wdNw7u+99/Px1Qol61Ab9ONLtlgf9dTWPK71ZMN0BkxxK7G0/TasDeBx3GRgV1QxlMperDcu
ivggau6YNlTtskBVOm3YN5oqdekiZh0VYUK8qCc2HKf6RE+roDqut+nBaNHFeGD2UEGXe3ukiKIU
8H0icDjD7iOujAgmuifRv4nOT/9juEr3aFGH3yYYHb57MWw35eZf0ItEMDX3vNoukipO0+UYC0/x
yVHSLc8PwSd+Zd7ijeEyTZSlmqVWM5ZYP0XWlljn05IeZ7hSWbobtXQTZ+dvW4MWSLmemRuvI6OJ
GYtec9KjJ/iouhSORfUOXErwO5j9hlo9pESwdbAn1y0PZLnV9hubQOTT7XYASbVfrFj6s/L2oVjY
8s8/cUfAjeR7mqEFcc2/qcd81kOk9C3MvZikACJwwe+n33HUpr/ULMROwDotJ4rTt3t7FTV3SDyq
XzcRdya/O3EJ1Tis8AGtK7LPdbPMIT2zp6lAtMMs5EHyYuQhrO0zkcbCQspl/mp4fqlou9H8dyMO
iYbQ1+tVEiq9qmq/ag/YNwYZlDNR2p1PXjTMwJbSqkHpVfNzwrGOeP73xhHLWEmZO8KNE5EPqqp6
yNJ5RsYvpK4YC40BYuPF+/pas3Kq6b7NjEDdNgq7Rh2ViSeEplWjxf9Q6yByxV5bNILqXxBWA08V
vJPJWCrkjUlb44/kVQ0lgbegwwLWwmz9soAK7hxE5dHbzTxqs6CkmEvugarAlBsa7lK/ddbPMFXU
l1S9472x2C7lxJ5cC//tTmJ9HFWAqjhNP78Tw14UCflw123dgpDMpE2/mnLYBKXslOUKY+kGkd6A
+MbjJdHbuAYhMofqYiyGt3vhXNWE2yqtWweY9dD9v8IMf4fRxeYAbSNP45eZw2VZrISb02AK+NdC
rNsaeuJimwDfaeY6yv9lb828MGae3WJjgsfFVmoTJOMt0AAkbyl9BxmAwWNc+QeFgXI3V1fmv9zq
eVjXWf/4yhq7cXwPOK6dA6hSMdYGfYuR/II4VJXkz0r7h+wTXYLK/StdznSA/PF9mnidDHDq42Mf
KxtfMFQ/qRFVJSJqTNCTk0wee1uNLrqXruW3Vvtk40hdcsZsk6kFe2VIAJl/+dnE6VDf85uLmRvy
9mYn+2viYTngAlNNaJ+IXJjt/S7WxFZH4En2++OYfjH4IlVS6iyY09XFr5MWg1yeZYmELGgghkdp
rmjwdGk38aKNj/dEtw4MhRNAkFC/A4oP8U7CjkSwWQ5uIzKwEh/Ip+TRdXZp2p7GaeyLtdJSZTuo
remsaPyES9X7aTGc0rwjG6arOzBo7GOn1ZY++l+1wiplGL0j/HOoxJIrsZYMY4XcmTGNwunxUiPy
DgwphNdnR1oE1nKtWO2KMVJXCJpJw565WKim98IghvcABhukv5uuQ3tv/vtLKzdkTih9ayVgfyxf
6Apl+4HjhEcDs/UkydLshpZWLTTaGFNDFE5E+naMdUiOEsQD6N2PmPcxz2VrT0+qbbTtzEkB0GBi
eIz1WJsogQeq3YWPAplr/BZAVGoa2cRyvI7cGarGKsZqw8EN9gNyNsUVlgvHpZtNoW4QVayAF2lY
AAb/hKy3N2i/aFWuLSMNZSeaZPxNPy4mRDnIjE5GBppp0RVTiSMmrYAFsZMVhk0pOqm64a6zLnFI
q/NME3+JKGXqQTAkNoD6DphupMzDHXpuQ5oi2nR17u6VHlM11C7sPv4reoOW5AZxEasBeDjoxwNb
BRBZw/LCgE1aayw3rJfnrcKrY6LzQfpHT60Qa2Vyb1ezRVAMZhH22jvx9/3/pA4hhtELS3As8LPJ
I0gPTx4kWS9uGs+17ILn6eVtWWTMYMaB3fI+95AIyGWQTvYItSZN68+ri45isa2RpepgVhARMJ4W
ThRnw/l+WghCRRxfR2eIuGMpxuxoX0+UzQxP9JfFeGbexYz0SIEPz/67JewcwWU9q5f7Ge871Sxu
vKeryhQb5/uMQSb9qO2otYFxAIILMIRANsQKuK/vIrdaLfyMGr5niSZeJBUH6drsO8bnm5Siza6U
ja9JhV8rG00l6NGyYhjYzerpE+COJXTBMzG92/8mcLV0Zt/EQkOjy7JQFFdA9yuHdnxCSBAQ3uov
CytJ7WTgBaM+QgUqlHVRiOQvbcU0fUZudYJldkrRU33fIw7C9RuHDUZkpuk2en/nvrhd7KiqnyJY
Hk4xXdQ7UMFbMTHh09i68dbH0C4WjOeEhhfL/LpRBDRcUZsabaGltC0VWIThDMfW4eO3H2dXyWV8
WRc8qpfpBEDQ9od/XrRp2ddxyedQyB5eF4jc8yeB2qUV1JO1Gf8b+Z5va+xtX/zuEhPaGdnLuUIH
AGAWWrURBAVgYabLf1e8LDoIJ1BzjxLw2hTYkXiOs8sX28yTr96KzX1FnDzbiKj8PAjnUIPvfE8C
NcQ35tRfQEUfiPfvecJqovy6Q6/5FfrYC3m3DuwjvloVpG4QnI7PjDr8Ka5fd8THk/OVjVJpEvur
r4dNb9RPx2IxcXfXaZwM7DovNm49vQHOmdCpoB9Pt/IlGyzUHR3wllU4N1ZTvRi60TmBj2vW5W7R
8CCwTYmJfXvXz13VahVUvBy8WCADqZQaOBq0EXsPW3cWz/9WoaHhMak3FCkr24rRL43Dk4qab3c3
ubKSz2IsvFLsgUsNpWncej+cC1GWRS+K3kKh/GX+6RhsfHo1yvjMS2k7GMURg3uEj8vGy099JMFZ
54u75gwNydm2FJzUm93HUY5PGl8WRGk7PLZzohA+8/kBV7X5VrEWuR3mxsi1dh7Fm34fvDMcyzcV
JLXVf3xqxK85YkoP23++akJAJ55yoiXvvl+S5ktzM0vPnIaP37c1g6fO30P8vSdCP5v4MT6fGQ14
DcEgb/mdu9o5efTVn8r9qYGTaM5WNPYf9uDIHKnTB3Mi6CuizTJYUSNqhEoIf4odjU6MJhR6RMAJ
rUg3CZDyAuqjW8CTGjxvEAb3FK1oKrO3s0tYcH6LdyFxuy/5u1l6bABhM2WRyWZIeS66DzQFPOE7
zNlyzA5Qjj2fRXxlTKgEH6VcC8Kbai6hvENta95FP9ikq7vH11TxNwXdt3MrJTu9LOldgaPILVKb
XRcYFACs1VGEZXCXWOknqFCT28HFrgsx9Ur4OYXCE+LWsj9T54luwfshYQNsZYTIRHDkbXpJJR/c
JZuzn/Edr7OU6xPGvrpLbMX59wqAxJweJE+0FhauGsDdKsau6EdextbAOb2s3/rF9sG77pgematk
wB1vos7FivImP/mOz361IY6fKcN1LsXLLgRG+MFsJ2eSz32OeoqXDThkCvq9YVaCGuHuxbjHn/T2
J4PuyHUmu/WdTNu5xbhmsG58e4XGroUOYfsEAc0zJwJwJkuL91JSpEcoDV67oE2D2/m7JhdG2FiI
09NpBPi+e+OMkXJedJusuFVuCFnvenV4mZJuv6rENdC4k5lb15Ddp57uyKpm9ruA6MygkK7tGPaF
/yoixa4V6N0uIc7V32/ytvcscgSsP1Qoh9ZG7xibZVYii5MesQ31q3f7Bn6ILg7Y15phqVXzFhax
ruZ/7crsk4SL4/kWa4U4k3yyprJTyKx2mQuQOo3Zz1/RCR27c7ZcULVkfxgMveTgL8EshQ5N9S1J
QLeEIRwsSKne83FqgXxC+7opH2gtSkycnUUVdawvqOFA6xQ1dIk7CFvCp92VHeswYjD3UTZne93A
I530k1ICYgccGSVvubO27jsFBdTwoZ4Ui9+6nsT7nlRsJg/bOSBYQd5SCIxByNVcorqZM0/X2RGr
HWck2cbIPdTLhVtF9e5tVhCCsa8gbrfJvN15fuFRyr7cgHAREzuSXbJoYDAPqT6WZl/e8Rn+U/3c
XX+ZH6ZF//6KP+4qelQ4L7iZpEaK7KjkvsJ3g7mlizZrtMoBH+kMr+AgMjaDrILYGW5HpoSADXVS
yW8B1UaYzUhTWIwAhZM48GAbuf9E9J7yv7sjjs2UxJz0a0og+wLd+5G6bUp/ehJjiBhSOG77eG/9
cexS49ApYz8NwpOcMqifHYTlXo+wT95Ajpq28wu8hiCNOF1bHBWmrD3tOQZYB6BKT2jkzNZmcj2M
n3K5GrIz84JGdYgxYIxcoblYh8uD9jb4nAZJQMdMdRAL0379MP+ZMh01xGeKvsdCMQxis1l3Vqby
nT2PRBnB2ETS8gsxpDaNYZAfB9TcNYwwkerQC9Yn1OWuZ9ibOKTzndTqB7V1OvbhcbPTwXWH+T3V
L3C9n5An2U+rI0n/l5FCFWtMqqRFMke+cSdT8LhWH4KnSLIg6GhaRblGSW62hj+lYmBYily1q7hM
dmFaNH43Hcia17ZVTkMJf1R4dQ+/XUoRP0PU/I7a7Q1K3TYPxXXlTT/IChDiMfULePPrC+Idivjt
YKDGJu7Tf7XpAHRmNtoSFB+kAKPXam+ggoPLHrN7IPm3bZyfRDxPMDZrF60H5uxLsmiMuLWYmlwK
q3ZUXPTVTv+NAV0X8lFGi+nlh6saz3i43OHg7HIX5hr69nSQz7FHf54ZETinAqhw5rVblCp4lb9M
SawSEogIgZAauy8dDxM/qNNhVwaJmM16YBOcU/i9B53CBt8HtuIx/Df7dgB5oCyPx2+pUHmeinyj
gYNQmcJgmeQkbYs7/Fnen5wMQkZhjBKVEKgKo/4dcQ7p5QsW4FBmdnPyMAhGk8WpR3GL2ujPdyHB
cdLy+LCwU8koKVvdj/2QNbfAHsmY2KtO5aaKYPC5PJQTSmtqbimL9iMJmPdSdTwccQMs6fgrTsLq
dkIRtMKs1ixW07FOLjVgKQaF71wtCuwILJGPCeRhgVIcE2q6MtwYmXLnrrEEGty2RnjNjWUdP5Ev
qdhMQQ+LRwsQlkkia//CVxEqUJSbDCPHaBX7QUrqszxF0Bc505lzfInLxa2GBNk6yjFTFJwfYWPi
fxhw1KHKiah5xA0MdpKOs9Xsi+PoF9CcYotlcLSkSjTJOGb75nADpLVCm/IQDgEd3DJoyd9caPOT
gE6/fAUOFNuXJgg7Kc6uBkx0HjBVN0iMCoxVx+bDb+h6LnUYg+qGEFA08fV+DFzEy24PyCZbl3fA
C7xp+RQ9MeECAOdRVRjOsPuNJF3Y5wR7yDF6MQZHou7BovvkYnC1GelvuHMahnqivIrpk5RiJuQA
DOQuUMON8LIE70CQQmETkV6XnU9ZtgSwB+DH/xMxsmTiU2AjlFYwRWSZ41A39Ee4VBfWv9oQCEg1
qZjAoBikECBFGhu2w0mgik0j6COfFsxORpDNx9K92jNxTi0+XkruzZFvuUXNjM1QuKgJscdBuq+s
Ie6OcMasyQk3TZGCPTDVSnLDD6NSU5NJaMmpLBZw3Moyhttdwqp4kb0oHG+ydh6AtxYLGobE4Kw2
lt1XdEYEGsxRx2ZQLlJYiuyMo1VQ2OfEhITRmkQZ95KmgpAtsy1VRxPvzPMBJo1+U7ZkkuTST/fg
GU842jHUmxOEARtfmJfG4ouZXSckMc/pXy8LrPT+15FCkwBQ8utgClROf+C57YK8nVgZ8UDV5RDh
JBxXyGJQdvWgxQyKl1msp2y5aYUfufkMtYHPiCeya3LqfmAvspbIx3Xb7D61U8rPQBNSvHP3CUy3
O2TKtpJ/eknmxn1VDwZ+GFiqdH6Z4BS0fWz0ZeLvFHP9xhVG+WczMWtw3lXcghf8MzqR+1le57mv
8iuMjLjEAx4ermQ2CNE2JMl8azDlfbDLJVS4jnGqfOxkuIROieK/kxOA1RhOsyrvs9h9k+60+v9I
gnXden1WCR0dJeTR0HWymNFaozsG/+r1Xmq/zDrjJVXN896pnvZHUAGuNrwPvtlPPPCI+V2pkvsx
GAjdi+LGVJp0gmW7PbngwAKMl+nRgxaOeAhiDe0vqjKbVHI0Fh/MQOytsv7GZVpE4xQsSPU4AHp6
/JoEyK3JwDbMOS9QxCW2dKUGX+3bPTwEkyvjnV8m/jgKc8mg0xszqP2DUP6+nasOd81CtzjA9a9w
8CBax0usuhR0Jtoz0PaizGATr4nIq14m1kOQ21oUAm3xzbBPZTtBTkj7PoYVNSk2/e0Kwq9QtwaP
MoLjsOM0LZ5iOBc/nDaVeKHVYlk6JWenOAdF3aJujJFXaUkZ7bWXLtYhuxO5AGfzKQhXQHuWq5xl
vmjhlMXrRKa8oXrKChqx/xlBPeBXUNXAZfNFQ6sygbwrF+RASz+wA3TJ6B/f1vWMRZwskDB9QXzx
9bQcOg33gL1i46ek7zkJczPrnY8AvDbHzooU0OzpgzbLNlyg+szuC5SxYISi/DRYNoBnXiA3dGjB
1C+Gz97+KkAV1SaL8P052LAOyzapMMwGtMmT7qyPjD6l2ID3EKpuKCVnKfIdygTpXF8d/ZGQ4CSb
lzSKk/dREhsqyeeQFOxGGfVgXdJA19ygdrW8qHP4DnqSJa9dGA0DRTYFNpSsLRAUkBcUq81/X9y4
9/h4fWcIQTrpitCTDDgGd2haxxahlXSVocac74lfnfmNWWfNOCz2f6fTMPKBAPF6PWOXA4Zz8g46
0Mi9LJ/T/UhqkF8sl+E6MsMzs7aBjbdKFvQj4cQ3rCe5rc8Qmq14xdXpY1uRBNZ9lTW95P0t7eCB
7sEeMRloNfHj4Qdk53DftpDVPohDQDRUJchJkyvbeSlrqxqAdShIgbXh1YcuYH8p1L2CtEWiaYbV
nPcnC+2yd+L7QPL17cXxLu8lcocYfolY7lToCkyW3+NuSGJZNPs+2Jo4fA+3o1TIgMpo/xZYIfms
asWBtWdQ0WmahbN84v96hr7S9uxXKxG5QZJMz1PsdAR1+7ylmvqeHBu9kj0X5ADGARJ9Hwqr1v70
ZqHTXc+woo5YbDZPNLodw73E4MzP37il7MeGjndGu1Z9dNsJaWsCj4Rq8QS9N8B8uvOvAUkzwdgY
p8wMinWZBbbDDsFlFUIFfMexYehL/ysau/o3qvp9BqUQQt7T5aGuDzHoV4Zd2Sh2smjazv11QRZr
KVdquNx8zcGG/rtopuWZHUpxmyJAhPngwoDHCR34cKlqlZXdlJ02ZpDyuEhJfYWSasKn2JGan04q
N981act+KLiB+fkRVbiySqnqEEMgL20JaxtGrl9NGwIAVnbt4DlJY4ET3LZaQPQE1cv4TER2EmLj
X5DeB5TgGyEVoxHN0NoP0do/FGSYSFSwGFno4MJK+9RbIqoZDOYqVQ1B8Gq792Z2b/yHrQ1B+Ruk
aPPkmwjCVX+jBJiQHCSLp/d5YXEmCcO9bXWv22ldAqTOnZUs7aNFNNhO/vMPZ8+uAqA3ArhgKqM1
aBVeSf37QNaiTaJs+22U23wQlrlV8qZj6noNKhfaenLnlmuZHvK/dR0jWl1Yb3ssWx3al8QtkSBP
QBS91XX6g9aR2N/Ctg6c7/7Gb2IlwCLdKPbi318pId4Mcs7yz0iy/Rs5RTacDx0WL5f4wVPtNKpv
u49nyT4XmxjspDjYPpAtBm+g7X813rYbgGGB/1GwbjUrBF9rp+pEKJHzckvduMjFHMQrOo8CnoET
NCSf8J/sWP3blSMKslv6v/gOyvutWwgyKJYtZxj+SY0v2FBQmcuMzaslNyYVRWzt8mlWWa1jY/u8
L2Sv23MfNJgEbwkiOQkUt9RBVFl6mGzjxJZ6yGZeuFsbnKPPjNrfi5LH00rB2nC0tiS+mam/J1Hu
a0K85RinlKTZ6OIhrfpiNyjBjK6j/RbRCUS5o/82EdmENXZFgBFs/0+SJrs9RofC3IA/ArnHjUp6
c37vrv5TY5TluMI4g9Xw4l+3HFsMidZrtue6o55bitbKZdGCAmUBkeChIsxQmMNnMPGpVfvLwZZq
xaAg25eucjQKEg4smnzySjubDK/bVs6Y8bewXPia8gwyvXlBBfUCD4U4z5SOmDTV6YkMDXK6NNlK
rXrqg8yZmYjQLYtcoHqBZgZkNmMV+cKPCpB3BZTTL3Ml9gWdOqgfyaDQZiOD4oZ2AW/qmlJAKhMd
fEkXQXwdZpmhz3i4qnNhip4HAtDSDK9ndYIsvbQYgd+k5TGLKGX1J4T0/P1pU15IGtcTlfxXRyQK
llP7nXcBdqhDYBQ70f8iGooVIMmdBt+9wY/IDgrIZMi0pT5/HPFoESz3dYIVbiJKvsEobLTR6D7t
uiIortEahWXyuZFAjfNvRzsqAnqkdrDzPZN7xuC07O7vqIn+prH07JhTTs09nhUWEEfvKGeebijb
djvuwdzgAx/oDDLwr23zs7fF+ykCNaXeDEYh7kPrKX4Aw6xoTKW6MwsXsF69WrxZaW/50Sat7T9M
38YJ6wEKKbN3kQuYX5Hf7F8XhUTDjNr0vTb0Q2oVK1+mw91DYiH0kE87k5mfhN6YQajbzjW/Sh5/
Y3sdi/3z6t9DFTZko19kF/pDMlrr98Nf6uPqyvGKAcRRC7AHDAJmiq5q44sTUnCOV43eT+K908v9
VYNy2KtbLDtSuOVav9r/yGzDtv03tdzUVf++EaXqIwksCqsrNpP4ZXLxl6EEMCfg7cIk+WRV98Uk
U5ijMVf0f2pOKTyNJskwmTpHwWfwmY1GAN2IalkuTPh1FUWoYbHtgGYk0gfhfTSoRo6L+0XiM4v9
EZgycOzZ5ipb4w3Vs4BYglWXUu7U5iSMBQHmsjQBmoDjKaEm7Stg2Kx1goBZ9xUb9aC1vE+RdV6T
0wxqaSQlDhhOmQf1ubNpb+KHLSNvpAOJlrbqKA+ZnPg88vgumdSUNdaBPVjm6nraBR5DI6sjqI+b
3k3hKo0Qbc1AJbg/tqhbDiIuvnr24Tph/Krm1/IcV+mu9jIX15k3RIpQCKKpmwb1pzzT0y+OTfd1
jCTf39Mj6W2LTJlskfuFzR9I/yWVnGVcjzhk4hcUupPoBqiULJnAkBPGckhlWqPlt/I2nLDJ7IAq
B/MDk6lGmpDL1DR1wHx/TT5/Y9ZREPRNaB/I24YNzQ9mXVezITUFLVe9QfyVSrzniWMzghrZtszB
tGGXhYKBayfK6ZX6RQyMMoMfUwz8ZXe9G4pkLrrF5Or4vfXVQ/56oHNZhELcoYuYpuKhOQNi9Dcj
Gp/x54fJIBODq+0aiOScoKO1dbtzDXxmJsLoPs2KRbYExUHBEFH3JooW22dXNIUGLsecuLDBTF8I
1A/9nJoPbveQMc7wdKwtzhkEUmUf78bLQl0TURzpWflLTo6ekapWHuX/wI/ui/1CoAqeZ7gY/zy4
v18S+x/Rtp2jW141Bsc5PBVER7/LZW5rqk2ShWyJjbh++aiErIjhX3Kt3/61UUYIZ4hNTjjqOg6X
r/UCkoZ1sFcCuk42Hlb7aSVP3ki4kLT420Etywk+mClmR8PKiICNJSTQMEoNqogIwMxNdoO7BXVw
PH+JoVIU2PK504FCfhkP2d0v6xYeMxAX7wwk5+LdoSVuW0x87dSbob7ikDq8gk2T1hFpz5io6IAf
NqjP4PXUnqzcayOQvNDPrTj3Pc1KBA0BEVhGdscteCsFhGtxSiqx3sDLwj6ejh+dUqI1c4w0UbyS
0660m2RZBlbis1VmHav/VwtM7iyu/OVNKlkmcaWY+3v1Vy7ISQo7m7WUIVvlxWVSPTqzQmjIleXA
dPqQ5tWuTP2h8z/7ynzxfENTshhKmlN7Awk4ixbrT+xaxSD4QUryHpni16DdYjyQ9xG6+oe1rqCz
tS08GTOml0s+Us2EAN+P3i8kcyxAhWsnfgjrtOzrvTYuwOJEjBDnITwr8i3UI+82+biILADT6xi1
hFoWqupe2BqkiBCxRyP7PERDBuiB1za9+aJ1eVam9gPGq9oM89EaHjCVrzcz3LaUkqpQaKcFru23
YKeFIkLzFeyjjjoLj3L6kSM1b/Idsyay1PyGyvESYWw28PanqZsGX2dVNYeV+pW49ED28Bfmjiu6
LPQzXI8hgFeeN1fuM8RCsQV7jWi9xY05bv7/MRNX9wB3SosJm+J/h4HceuH2e6c8tBjWgJ9LDhrY
houbzk033vZ8x94UDDeAcXorkpNwQxymUnDMwwHARk02JyPlRpHICpNmcprvQugMJjHBjESoPq4U
FkCFyTC1VlMQPBdMPijP6+HCDJuq9RyhuijbMTg1+0mDi9tuwuOxmqFSCBftTMQTbZBJl7KkZP+/
4WdTkVSRsVIKKHo/VMrNOSRcHHFuA3C3FwPwa8G2jTfhwvwQloB3kyMzBZNpsb56CIUITcXtQdCf
oqs2kWCVLKO7Fc6LN3xIwc8CASAhNApi6sjkKwYCHxZX6/LqEpieXBOuW2gwZMDT0wxbcwPST321
YoQMVl51RX7bYEpjVzFIYaNubw+p4X1/RyBF0dVRL2bOSZ98rlsw/3fmX8TV+LSblEo792sW/Fyo
ATIKrNIfGF+/mB6HRkMILn2rlX2E/QTdhyID7hFsWfoqm3wAttDoWj0BTcW8GINZPwYr1yXk6Fjl
IzvyOrtw1VpaDuSok6Qd3pTVCC1aLIAIfX/x0F4XpyicfEKTwUBIxvGWINmbhc7gYBciWm9IZmU4
zShHzUzwMEHSasOeJfHkAvwhpp7Zu87yUO5VWIq/h8MOhpBVdsq3xAZeST70q27+VnQ3otT/QHEc
dn5qqoG/8nkbzVipEpHtCCqYWho8NsKnV2NbL1KnNDvVqwRQ7c/MhC8o2Xn7iEX/IJRyLkPMfoDd
Cd5CCMb24OlufEYvtizsz/onhE0FhMuJs59GjnqC8r1KwwssTJA67UmD61jG8i+WFaLa017m2hxd
4m09RFz80uXMTPANun73ruzjd1HvAMTCI+kwprd33T774swsAjRFjkRegms4O+6N/mmbi+z+/a6S
82cmdXlDQoPueYeKkdQto1uxZJ2ZtkwlUU9pLPXl4XEOtnGvBxm09gYcmsp1Og9LhZOJYOLJ21bE
4LUm4tV8sawv4Tq6ZXaEF56HRXF3IoHquv9qskGacTO8WD486DAijAmd27FKUXiI9tqfLtQL16HM
dyE0nHJZyGlJZ3JqHcLWGcTvW5aBAdj9+OFuTnd6S5g1qcMYE0W9Knt/flh6CTTaptA7Opz+R1NC
hIrh7e7WpvVDenroYITV1cOew404xqT3Dj9Bwn4Se+xOK7XghYC2IwllrZyOT0swqm/l9eEW18Pw
yGLPnuBmfL8O/SwzvDheLtY+mrza31atfdmSPQkLiz0+eX6J79Rt75Z7hZ1xLaVa7P/Ws0cJGUxv
HhzdgVyEV4XF5ZoP+ExaKgLBMyaUVJVXzWTavQ0/pi8juIOwq/GBZr43AYuFGLojpSmhHirMBHER
nU5lzDzQIY6p5I3e8hlyeWKghtQL/YD/AzMTnzMz/4YnVOIUR8w6XM+tRE2Eg8b2qGmMRO0a2D3+
lTnP2oRP8/aAs7Nvt2SOyjgctUXKg2v2VHQLrcX1HXvIFUXC2R7nFulRDjg+XgyCpl70C+U9UEii
NOpo6+7hQ3PT3qqjMcDaxNKkxVmWPNkq5wlqG28K52COEnzToYqsVEOSwYM4vXKhjt3y8e2IV2X3
cwsT0sJIXX5iVC3TKqpE6s9gz1YRe0dM7rQzjtMyMHew84RDKx2whHZ1t0MrjhPqU6/yaX+BtOV6
2xSCPGCzeiwA1R6onp/OOERIuuuHiN0Zuj7MG6ToXvrkuCscR3sg0iVrzyktHxn3/rO712m/U9O8
QZ20zna3iO7Nz+5ATlOvIFik/BPw4QTW7GVZ6cS4ezuIf4Ivbz0i+nz8Letl0VCotzwpiJZSOvWN
wq6tLYEHkkNmIFQkasSuOjwq2bN/4fj1AT0qCxqEGzaZjrhDBNhWSsU1u4BAf3IqriXJ8i1uDY3H
Rk2/vtI9T8vttYRe+Uij5z+5yJzMpuwde4LM8FUk+zXslNNOWxU6XS0R+hTDR1dJlSLtp0rS2MeI
wX6+M8pn8Ov2lloW9i4HlpWZpWXG+CDveEflbmfzx5Vl2zXxK5ShFjudJNUBi5P1DdlKSf8/UIic
F1heHUgHkk+YXZ/g/BIG1dK3PXQT0v1Z+Dl8kjWLkyVsgAllAww8QsFdmqY/2dgdff5rLMdCwbXA
lV1y9oK5rxaBADoOLRLVmqWXXpPAK4NDTXzaIKI2rZ8eVt3Jfkm9LHSEdfGwblqTP9AZYrPBxfUb
d0s+6g55nVNEgZ99CJqxULwKAlCUVPDwYCWKH/i/L8JhOTFGfdNHOB9zA869IpFqdy09tvcx20ZV
OPIf16aN+an0nHXcNVZoXk7wCVjreEUD47euCqdx++OQeHGyeEcM1Ucfiuqxn4Q7W1bHWskYJdY/
xb5XMzt94Wt+xj6Uc29u2gsxAVNaH5UUqnr6KwDuHdYuql0gnrxnZ7Ulu/VNapx+OMvZLnyt1TvK
oRwC3l28P6jwhJQjpH8F6Bqdcrdrsn2M/wrGH73C+eBXcQ8VCehr0kqO3I2RED5VEy+ZXc5xD/7k
KZ3o4r+ZuldGcLDCeQLbzQOV8aBYrJHmZqQHj3/rqNHnu0MD/0khjqUSRAEWi39mh+JnhQD+S+P9
6ZGP7QYI13pC912kJM0cV3Ra0O6iROFgY9CIaVLN0xF4cJxyz68H7Kdx3sEHMdOBpbgOdgIb5dEC
ZFCtTnevd6t6PtGJjljoN5Ty6bt1CTGKiPQv0QZnjyUk65cVnRVKKfk3ZXaqa3bZvoWtoxkT0CAx
pFbAHdDZxx06HaY73I4eQ7FI5yYvjk4RyALk/+Q304xvbCDX5Jm0/Rn/GR+/h4NSiJQDRQVwCo+B
LtKiSrnB36wmDfpWpxcfDNBTGfKjbJ9CzkOiyLEXKjJNov5uEfl67y0nczBO/Ayk+L8O1vAphxMm
16AJqdSa3J04Ma/EJ2+39QF54D/Sc83y6HRak8pMCQfiAtptSJNN24LMWLLGkHSkdWyBkArXGQnH
0qShh/bBRNitjSeQU84JCnQxQkZKrdORDrtvGKYHlh3zAxSNmpw+LILrKwr2lRqWFNvLe72yhLCp
pvJTaI09P4ZfgPrf2NfNglJx1Fl51IUWC1M5ByqX5agLAdiTtO8omo/eEakcxhw8JgHyTEjFAlkb
1dwTmaUteJyN4F3nEooXD5XShsxc/URWhdUaqyR4cvvWZTUxNV/HaWtWY6YgiiGwogJyv8Zy9WlT
TIJ9diCBuz1/56pMji4AjdzgXwxW+d332LLsPmjRYnUV0wS0Mlu/2RaKMAlhHDKhZJTs3S88+LO0
odO3ejfIsULD3KsXHgZy9+Hao0FDi028ra3m5wvipNKn6wzm72bvpNwOeNLM6x/HhUqRLG0culCd
u2jbbUjtkfjUCSMHXsjrqjqTXDITHA/tI6R3PF56IfmWA7UUx1XrX2KJZxE1kBLrKOEIx5dHpaiF
DnrUUCNTSJEivsvVXfWZxrLnGeCVhGokpfOXXkUBbEpyHpygRUggrWCxAX/mer6jO7EYwyT68xpk
/PzmaIWXrXADSiNX5fl37gZv++y/LfQAoyxcRrI1tzNwoxKoWrd3aLi9wp9tHicby5hlwkCdrVsA
BP9agTjWtxdR5dmgU4eku5j4+F+kluMeYmGV8en8gZMChCV+gFGRNiF1bhnXsqzB51Fc2km+cgVy
02XrInwya9UQWh1bDt7tbl0KfUbv7rPuOdUGAK0eXPmVC/iW61eSk9SkbSKKw9N6lJYfePiFXVX7
wTvlq1KZwfCAroNCVPZiz+xejRQF5ydgg11/NkBhMDlsCy/vBgU2n1WJhTWH3RNhhL8s0NR3Yv1F
jNli0osZ+5dDvndyTaRpGb+WSWXBhHm9BQoNZf52Rkj6dfsxA2ImEjyKXrLZHWj0o3buGAs34cpj
plIayDH8VTBftSTaGnHCdRt6cciYFiwRU9cp6UyAQdlurJ9zzaop/dxOOtD8OFPI/3lg1vlcSGyy
4HUVY6nL4xncFg3PenqcI+kNXmDKM9FROO9whZkRpoAtNpiqlwRQO29fRUhDSF1p5CTdfw26lEtF
kYX0p8he8kKX7H/6lf0cC7WWlkbYlc23F/vAviyJoT20xRVQ3BvmXVBP7k76NucOMt0kj4eYJrdL
yP2MoPTt30qkTKAcxn7s42dQA9j5w9FLeKez798+7ouYmMzs4IqD1xuiQif7+MSxtno2/LfKAo73
RHHIaO0RUAic8efdjQc+8uK+rC004U9/yefePAzGtalhBPOCisE75d8RntRkVh90snUUX/LswSZQ
c9sLNh7Xnx2pXSqcVCs+r5GEYMjvU43SPb5fB5JZ/2FEB8+CmD6+tZDdbwm4C60CRnBqiVlQMBB/
W11pC8EoNjASV8g+f5k5h0mgbkSKuX/WhCK3bc6DxJb7xivJpDJG/U19cKTj29f2MoY6JJ90MTiz
5ATc7suE+IZ+jcFHTLZRjOXOiS392hOpIRoFblwIeoM1XhhM8DBjleeqLL/SuNNh2xUTTFW70DaJ
vKWX3bmQDoJ32HYXGonTUrRgJwAJI+WW8dtycsy4AKuNx/0tD9a25SXXWQYvf7286xiDUgF1Efhl
OJTMIna7FibfBOppwEknPOBGVVtiJlmiT1yHHooIZJRpZvARs14K1boU14bptA41/4e1NFZ8Iee1
OFDYtcyBekkUrPhxI90jdCXj84GsjVwqnCJPG7HG1wkctHg19A70KG6U/PJuEWE0KO67lXodcL1y
4VgbM2bTLcQLWukOXBYCdM0mWgsGRrxicvJec41s6jagaE5UUqySg2ngCIixo1bXc4O0KFAAraSS
qMYZ8/xXsoIiMfu8BKkAozAmbmLUkU67EOkdF7umR5B5ZIZrVLZm+nQ4YZMhuCsqpP54emH5G9JA
KzlGqk9euNoAUH5h3BxMULGktkjGdlTQT+m9E9swE1hgcIw9Rd3dB030slgIJTILltnS6rveBbPE
cMNx43Fafte1gwXMolqkRrcZcgaX7IhiY9kyJxDAPvyQJ7yajjSkby9yR3eW3PsYq8ccT/4/WyyK
63wtDsBVac4ZAHhPPJ2It49HRlduuipI8RjThDl/Dlaoh1DT33G1efowCIHMGSb8jGCXb4WZLi6/
TY4dvCX2T7kULDo6Y28L/wJstvhDa7eUknZTsvnCQe5sYtTbCJeMORAq0op7MIiibWgdSMHdPWU2
0eDF8fmeyqCF5kCNjTkjc8bnw4CvmXgLSKE1VDlvaG85ZrLFOhd55fK/MUyX1qAXYmouzDU3rNqF
93v16LY4o1ZHUbGmxcmE22yUP3QkMN7p9NRyExgeRHOgsmRKwdn5tmKyIHq6KPjW8NRm5d0WEnBC
+GUP3Dr+BkeDFIelJPv8YM0+Hr0xjrUn9SwHDKwGjgxYaxOVxmztxmKdmnLm3LwA5G/sLCbbP4+i
TRLuu+U3M4G8ufsSk1ZdSp9P26cy2X5HUNJiqYZdhwB7l4mAwc6caUybaDewX+9WyBtyJwj7ySjY
rw5LJqMlaucsiX+Pwe/zWO/+jkXHssDOqirqsl+mLsdLsl50fuEseLB0KABBbWloyd7C3Vbqdrjd
DIUXfdueqewmlqS8ozkR1jljGV2xVGxF823y0GIXg439fFy6yXM+0KSDWgLxwk/huYRJQd/m66Ve
vdRZChqzhm2fYa0vcW3scOf8dvOO5uODUBwzdxnvzGfd67REeIG24fC7jYoHQlM0xB/KkqHfKW1j
qKWBS+KUh/XPaVdH0WylMA8RPA9pStdovF81IAeYoIuouM8EQl6ecVmtIVZw7O6s0SCg/G2m61w4
6AVFv1cyka0v1uPySE/HhMNLEo2c6xL2rJWTdoINRjxmXgovog0MD3JQs1VXsqEW+XJ0Ix5elDbl
K6dy0wi+3aFfMYD/DFCDqGZQZFNikipb9RZHXPKA1cKvDbuQi6ZfulIowdGd+UWAm8MS0jsK0L1O
Os2u4ymH6IKiBRtLb3eJ6CQ6Es6yeL96n335ZEpfA80BeDkHi6RMcKiU68xibUmJOWNWWt758dWV
DvbBjJTbK6VlmfRTkl0dHlRU/JyGdrolucxWb2yNlPrDDBP3PSLyEcawNNFVNkY7VPReAGl9LN5M
JWGuOB7OOJqf/nqwzD0eFSTBQYGiW+rYL1a223M1xO5dBWI5TYeJvP9YEhdmJG6pIPRqWTQC742w
J3qI4sahDcGx0hxJlvLPQJHiZUT83jSxNPh0CNAGyif7WUbWVnwdSvqHAac1lUvUkD5P2IXE2qyx
l8/+YMT4oxB2WloeV9wZWt+k98y58dL5RvuMld0yy2Q4JaB4dAP0M8dxgvEhC9PHZ8VTtjCQzZva
K0Wcf4aiiyoefSuW27tWFTjI2Al31uC7KyPbnT4IqjmN4HTvwFCAQbRDHKQAF+d1/S7Z9O7q3O4I
+JnYaV5JU0Wy7rdnU7aTNwh+cz2+w2Mv6o5x5TCIRLU+LEqHeNwYBZmI5PhgIQ9zSLrXn7W50753
H7z9xR5XdLf2bpR2C+j5kn8jnHtb21topm7OqxSz4jtfUuOXgbgveFhQHdwk1+hsKP6/uBsBB18O
i4UhvtgVz2WpSPVcZlzh7mciHzYNtqdsk0EBkxNaNzajYl9DYwgrrXuYQWHScAXhYJVjTwosyYsM
gKMLBmsxZTtcUucvc/8xzggfJcN6e5T6v/6SIy/UhSXWQo7S8ECU7sGYc63rHPf1i9CKMYbfhtHa
Vt4CeV2IH4Ed3lD3TwjEQZ1NuxaDtyj2R1DU2x8f+bNIxGT3yDCWUpLITSKjzYfdB/hJ1M1D0ktP
XedNMfy7cAQ4Y244g5CzXbLmslJSracDdr8m6Jhr6e6zatWapv7HQ6SGHV5IOkE0pfEYJaw/UNSO
WWQm2VpruEPsj5d0Scy8Vd+97BiTqNv6yY6QzYzTyRBXJp94NZEl0298nyleAQhmVRUZYTpWJxOE
OBkzW14zmTJ8heLL4kgEGbn9KhJoB+0IraWQpZEXPp81Nq3E/ihY3UFL39Uwrp/OyedNShYobJr0
Z/P1B39vopzw8TfGpq646qRYvqcKAGSyQyI4gp//CULsJsAz0LD3gNZ7pgS8T6tWvMjwWIGBfuuu
ojTBwItXf5itq5FRZzyWMQqrKl1SrhtUsNyEBTgSF3c1HoE1NzzTbskV24TpAr/uScYVujAczrUR
19VbIuhdFUKn+JPamEjXOdBj+QL1TOx0rPJRUk8pxwjutR63ZWz+J1rquLmEtM+CRgnVtxUASTZ3
UGgWtvQWhJPsm4bh7sEnSZKAfEx8435WHpywnnGN1mU9nyYxt7zUx64NRjBAb92Y7BDVUc4fCfsX
uLSunZyDjxQyoC4bo4MdjklnMZyPWPCm+FN9AiCDLQXM/DeAtDCErCMyJqtmTCGwMwUVIh3X4m+a
EyGcGzhwqAZpYt+NSCXvKSfHi4jPQA6oRBF+vxo3V2vR3oQTyaz/hZYUAE8di2QIm7FHmOS6Q65u
2kDYmer6OeIzRTNfQA/4HS+ZkSKNQS2fLK2JDTgPkdAIKaWUqTo7wAPdQVz4uXFqKKcN210RnD0k
K+BX8UJ1GzV32HJecEM4QWmkittrtyWdesgFYc7VidZwvcZmvDvzx114/xq6UOvc5+zD5g2NHlte
MkKGlH7sgkOhSER+niRCh4ImB/DlrZZCJ8ylE4KhyhaaInJnzNFk1wvDc35QuJQTK2QxWOckcwpI
rxbh2I/kFbBOzhwBrKq7DcsJf/2Mv4rnpWD16ZLFlJbPuOupJK03K7Zc1lVD0+kVnpAgTwdRuyqG
+QySOe6DX8dxzF2FQ7IR3v2tX4RkQTn6MAWfkyxuRczSk7TD8PHg8LI1o7qiVy4Ggdb/QbG0SQ5N
QlmwE2pOKt7JhGoTmrAq4/picag7SfhjC2g28lhoNHgLQWj5mQfHc07EUICJnsJKRAVNNtwFH5Rn
StEW+4aDl7dqRkHayVdK6WYKuedLHCT6XM1VLiLTyHoZnod+PjrGtTQNxpp+PbtWp5o9LoALA+SN
6nxW0ZnXL8j8AsnPzdEN9r7uAdP6wwFW/47738Gl9tFUZrkQE6Pg8TOU5/p5+JGLfqNuJnfAUvxO
2Ibav/Y9jINXjzRV9admE44JsXwB/zmPCST3Atjk0tEbfr8aaK54o5rkuZjSyrDXgZiXQSDyPV//
avAdfZBenr6358RGC1Bee9O/gERSrOQpSoxf7pFNZFeBvVf93ydkBz2sB/q2QxNgxc72QMgh2/38
xChy5xDrjswqV9vgpLYFPGvuFAzS8D2ORk2pQ5r828pjUzreYethywNvwkd4DcVtTTlqocPcTCXW
Z/t927aRp8OWYSLKbAiomzTc61ZAKMMfTXoWfL2NGrZuhUohpglCIxdM/n4o0OM2uwGnGnwNMeVZ
iUCBqxCY5F1TbVxi05BrFESxGX8xvFILLFktpUsKx8FeR/Bnaa95tMW24QEVI9yBNH9liUZv17Cs
EiR5eFSoFZ/nvhNh69Da/1CktHlR/OgXNDU2xRoidDlTUrZsyGZzA23yeH1PIJ1EgKucy2BRqE6A
xqTYtUii7Y+w9Ox9ZCV0O6rDzKcrWY+iZDIq3g679fhO4HcSbvEbIbD1WSCtJMJRIGWx8cyHkzwQ
xOqa/mL+MY69olPiICKliniy2i6UhLxD0hX0FHJqGdfoU6ID9ivsl/otUQ8Fvi5RiMmBJ6Q3Mt01
0LjZYgWTMCtbbUoMBG+H2kmkYwSi2FKj2GmNU0mLNxl5v196LxYiibWvFNyCgHN6HXgplyV+KQEU
coEDyxY8Vd9dElqz1503A2xb5BqjQjhneTK6XH7rbtfQRT2LnNRuVY+kvxXkqqRsst1Nix84eGhi
LvlfaCNylCevtlgyiO+31SbDJkA2Txx7K6NiCd2rgFbYKWp88KhnUZ4qoqLJL/cD1ycJJLaZ6aEe
WB02iZc66Sz/03a1PuL8nWvO+D+phe92KBuryAO0I4jsIpNsHSe3n3gyWwh69XfJjiom+hAUtKPP
RypJLIqYNmWWPP7QluDRKvz4eogeq4WmITIQjFkdRAoNBuNwMKzfrBqLBHrXMI5WEfbKqP0GMfDr
9l5YY84h4uH5xuXHLhviVkc81gJhfvxyWDTcLPD/mDPZxzncxM9SiTMcUJIcehXy2XTePidyl4du
542WK/HfB15CrF5G2c1Fp2IXDk2SIWUhHn0JvCPB3B8Jir7ImUbR1kiqWLt0AR9eNEQTu0L7kFDH
aGVJpo0b8Qd1Ivw2nuoRwSjetz3yVgh9Lj6NyIYDU6BOeryBgZNSva2VzIxPW1/iADGbfxcSu6Se
PCTRceOzP7hkaLYK/372fgH8+tJ9PIQBYVTN5A+ImSNSwwa0uR9ht2FZM4fxh6rXGQiu2MtVqO+k
The43ZlulsnjVTJMNVvYhJdLhKAAq1G+XSPReRELaSTrKXj1gLBUlHXn3sgPbVMrIdPL3wtjGEpb
FuUo2IQgTe5i/5u9GMYo2988Sv4tAesJq5lpaEh/la/ZIdPjndM7A7NX9E4G4B6dlQKPasC62Z1F
Lj/PxxKoUA0GT+tfJPyzRYVh00djT093EAWC+HHbIHLJ4AKC7fs24UlU0u0hNN+XEIHUVVezhNEg
Lr9F3lT7BK2BXCIOTTBot4s66eWIeDipSHUvLQw8N18MhGG1PmsKvI5uyf34sKf7dnoV8gp4uB3t
f4xSwJDHiFYPZqtXSv//kOk71DdzJoKJEs9SVj6cxa4Z0Ae/DiwSrHZSlUXVXjE7YjuWSNQJdo9F
Qf0CFpqtX5c1KxelyTxLzcJyZjy6vpl9nf2nJcQv4uKtYPFzAi/R0MyiJakArgw7DctpjZ4Kekl6
ZSHhcLXVRIXHkNYI19Vl6h7oJChPzNoyCCV/gwi+vFvTG9mZapRgl/KseYZLY+9IRUfVGHo0kYvq
OeeQSFaH7b9UzP8iAvm1+AU/0oE9VaKPneXsq43jyIxdlbrBsAsZCN1UBjo+9Arq9lMtpD2JCbCO
sH9K9/zAc2zBZtJVIVzuSvxrZrfDoV893zKIjBBtfghgArATdmwrdm8PkUodPPA0mt5YjDZkSz7H
bq6hJWpvw6uBaVJitmtG2DHyWbvCSgQqSEKjC61uJIyLUmG3PyWqKXCXNs5Bn1hvv9+ft0YoVQ+8
xBO4ckFj0pY/rPtFg0QnjgkrmGW+7QbdTilK8KWLF9PrteNGxqTF/3KoVGpEF8/jL+AAJ817N9nY
hfbqf2N2YzH+Xk+xOa0PbErzpog/0pz9guy79Z+dYN+wESSEi2htiZHvqVbOvRL3SEn3xdlpdNjy
wk6U1gsz4FviSGXX4d30MYOx1synbeQBi+vBZuKlIsDz/t59nU+/AQpvE9p85fYMz7MXQeWkmH/e
Q33kOvXg4PLhLuNd2koIM3Qncl397N4jxpGcrOAro76DfwQT06hU61gfGxrys4e9ZJpVZnhS2dU4
hWiy9XB/XmDlHH75G5ERyvvS58JPJxPT/pwif6iNHwLrd12j2EgoJtXuOEwav+pd6IyC3askqZGj
Z8OmmGhL26RE9a1jh4Xpcc90r2t31QjqmFkVCtkm7BJbB0VXYAv1Db6jpFrOrnBHk0CFA173796V
V/fksLG4TbyjpeOkrN3JDywEVuiyERE/W/G+7B1gcm6hAvg2nJzoa4fMv8vtApc/VXa51pSN6Skd
t1hrB49ze5Rc/pZtIDxqgGtK0SvCtpl/x3cbBp+IW+8KIDhDSD8CDxHSxRnrCKKQLfN3Q3HLZDUV
G/h8Smeo3bo4c1QGoLugnT3ecN4e2QqQ8Mv5JpRvXvVDe5H7Jl1nKnqRru2PkrXGPn3JitUcym5K
Gc9oMUybwoeqMjS69FtnWFoYYgfJ9/um4NUtKW8oDbzOnQu0sLS/gYxs+3ufN5sFX2VTWLYF+zEg
abiwzqVymyO2EGlI1mGjq9cCleGP/Do512uAWvvZ+/IjQQK64puDqevRjioWQ8LFlJrX0W2Kk41p
RaYMqrICmzNblLLxS+40AOY0LcGX+Qwrzf55A50GVWzfnMsdJEi0et3KXSYhx4Ftrpd0E+dLgiuB
cD9timBmjOxxiqYdBwjBrTXRyHOIiaQAnOgJHcm38IGkZ8awfF06L89jC4DVwQ6QBZz2slcXjFBQ
95jr7tOf9Y/Ra7AWKWtRM3AVjpDT0nHXLOW7gD7js6KDWzFyKB7PVc0VbUy9KAsoCgSjMsxNcz0B
hjzsEwRgGGZKpQIGoWhQaxN3BNlkFgxk8DzZpp+vFhbHPWIuoKl8buHqDwq69xvntsGYxW3sgKzu
OhJ+AU+hVXrGq/WvP0hcxEEECi3jn4jEVeziizprDSo6hwixNI8xSqcl6MK5eO7Y2hCg8jXI/i3G
Maravej/5Q8ShppffUoeBQmllr3brH7gucWhrMM+5xTQMHEtjVFFy2K8oBgNB9ZH89gyzlb1StHB
Uty5dMEpNTJ1ctr27y9LPdcihqyhdxz5q5EoKMhzMFuD27sVFZYExmCa9Vpuf1GEPFr9bKH0Wkei
bK1D4DgycO0AwDctgYAfQAHw/xPyeEnvhaawirNbaAwQ80xpBiPU0EoloC6y5Uh1q4SZu0j/R5/6
JVUbdR5B2KAdU2XrHTRwnGxJv/EubREQRfS9x4m0AqqkS41CBV2chtGa3V2MiueaFHi8okrxQAfG
E93DikWc8kCxHjgsSBfwiCOdH1yCsoo90lctPC6Dt04ju9tnom2ObSOurExO8we2TVloQj82gmMa
gNZS6v3liqyk0Ffi2Ik5FOTYkpbuc7ZeOwqm79DaHaRXHVzFVf33rWMQghoiedkj7WHb6qWjNome
jRHJ8jt3SOaGxwWWS9ayf+rSZ5Fcaw3zq22UuXrsHKWaS9VuLhtKG5sVNorZkFSzxQUSC774L8k/
e7w/scNap1zAmJD6jjDfxjLG4zNPiXaXhRnvV7uWq3YOGRBoGG2LNBYoPpkA7FZnfZD78x2nW69H
gRZLvxwMJ+WzZkh1BhLR1UMNj0hfAOoeVfQ4S5zCXSCWfIUA2jS44ZTQ/Zu+cWHKiT/9I76rMJUQ
QfjljTZ4E8M/MjF8JV28ZoCllii+A+9TZQEOD3g2cmaUV8Lsj++5813z66g5TbUbALEBghQtXuli
4ZVVkgFhM+qg7Y8StJAUX3ZysZa86lfoGIUtgTVk9QC2XmKH+iFQ5dzik2ZvxrACwTAZJLMJIsV5
Hq9iWKw5IEPpHI2LXcyLmBT9kTQd9Oi3bo6eI2UMbp/Sv8N6SBpDsUp7tLz4Jpkkg9w5l+4+N6+t
WRgT30rvUJoo1rtCV2pE5Gp09HcKyI3ZGMM/GycSvckju5/w86uEDmw33uMO27g+BkFLEdbiG7hA
piv3G62BzHqOq6/IVdX+SbGgNe+PLQYBMr9uPtRTckg5zPJFCoe0pOpMMHxJe7nhHHX6ragKx6aT
0MsnGdz6pI8U3hhX5UybHI95fSYg5F2aUv3z4o+VupTiVReqCDU/xIqGQ8jjlcVwwkJO3eILLTdT
QkvcEE605oGcrcFg/1GhPNBaZep3/mXnMY9S6U7wtH/t1T8Gjo6HuSmyhGYXfkHwgrOEW4Ic+jFX
ca3wu9wX7ZzZrKGhG5JdObWZZfp3JVR0kJ39KI1rGweVqBQM2eIqtswVyTdHnvtDWP+YpdtuxMXi
YqEqdcXdaJ05sRBdusnYMXJB3HXBWE1oVF4dU6llWNYuU0MbNcaDn4It5VollLrMDjZEJdsidctk
rYzyrIAUkPKrURZPQJZlrulmyXRutWY1jMrMWhv8uRzRrE655YMOuHKs5c6VN1/PE0tMWM3JA/aB
EYvkIiUwxA1PG3ak9ESHCEKJpdenyK1KALZBf4TqBptIxKQNUpaeVffffOMzXM29JN1i7E/4hU0f
4FibwccBRSRHiSkdzX5uChsQlsharqBhWrMIodCcxcQwL30Oy0pQ44Z3NVq6aSs0AE6EmXv6frbO
/p185kZiyIgK3geT5Qulo8oQU8d3vaE+1Mqv8JYCL6nlz/narzbdFgA9BXyvefzznCecjzs3yaas
sLhaDf9Alei52nmhc5jD/4rgJ7K90M5ldbZK2fg8BRPmqXBY3kD0jyjaJwLW9ybpuKzcS/5NT1eQ
VLT1JClEb4MEnHUDS1IE42wPCNHvQHOwbpJ1h7gh7gwpUUtsvJgIorjOfhkEdMmfHsaj/7Vbjxw4
9mSfE5E8I5WhTUBdHP4aJ0qCmrIaQE2Cayndhg4Cp5X2X5wXOeCaHzdIi4kRuhHRwae99fF/Mxl1
UURPpxijDhorG2LsBHsZuVC6iwhglHOiQT+ThEm3cVU9VyRnza6eDUSuPI/hiMEwYN3w3x6uPGym
F8OwbXcYbS++vumn6Xj2bz081fEIKyZ9PukSvP9iIs6CCf8o9juaSG9jxRc/l8DJEJG7wX2urrXj
4GifmF2iwUTaKNUhdNV5MoV/2Nqt2oXJZbVuYhwYAI5XrEgUyIcIzBYNbIDSimrVrOUpbdYjPOEk
ux/PSVKg/+366N7061x9amdQXEd07cZb/bafj/WnBWvw1QDUbyqmxilDbGwnBUDv7EaoZypYP1CX
YEks67uhEsjzR8uCVKW2kJ3olS1k3jJXQDkLC0YzHVzYcPSmeG9HMFLupzcYiECWGfYxvoi/+wZT
AzjidbMZypVKg8JyD1QKSYH678A/gY1Xq28T3gBCW1XF2iJM4ngJK6fHNAHkmqfQ9q+I36VbQpgh
ySB6oGWzvhGlZM3bUCaDz9lQpStQcqbpAwgCK3imtpoQq0zSfF2Tf05x2aqBez045q/0PVCbQXaE
Tb2vJhY6QO6AIzF4cQY0TZT6nS4+l7Tw9MuGIA7bAmodsAJ5nSLfftWG7S3RGEwmFNkWQKuVIsK4
LqdrJlDkjL/9slUTPh+9BLFnWcFLN2bQ5z6EUb+ZsJ+6sCrjE9Q9o2EmXwUPSWqTdaduhp13+pKu
9RpWszShAwWDpbD4Ui8MO0SWhD/njcZK9lYOEPYYGQtOc/5WCVdWQELjbrRn1QI4i7tDqMNHs6ED
RhORhTWPYqDSZS11O7ysXZzmyTGRTNcKU8U9e6JxSChe+t6SwsQrqm5W0vKO6ktV7bfkdmp0s2Ia
6/p0L+SjnvHYZxWhXCHHvLvdFyTQ1/Yzx4kxNmA6qexZ5Met+iI4mhsDBvzoRITjiXvn3ZAmtcz9
mRmCphsg8VdIB/XhYaXo6/jzLRDmZSy5VgDcR6wkIVykcDs9a4TyQnY4GqU40Xiitcq+XfPHFuzD
j2JxlYGeBN08NauQt/ZtRhaGAN8s6H9OOed4qoSx5nJ/R0CxwN+Atcfqo7WUeqV7o3iogbRRQZng
vABumLuZqYSBlYO/AxVl9NUG7rT58fVGQzDiUvXgiqh3CjpAvUNPy5idamxvuatATX5tS62MRy3c
7q5ApBKT7K4ue8PNw/ExqVEebC/LlFK2hCyVXjg+iWgjtksWuF6hCXl7z3ph2Q4H3cJ8ZjE4HKqC
W5L9YOH5pSPo26SpuWFBn+W8zPNhb1gbh5VMqE9ZPMPks3YtkzsOiFs1dcUuGqPReHnh4NK9F7Qu
kXr1uBzIH88h/SjIweolsCyIX6Z6q5acZalS41qePLnxe2hxDuVthn72/nVrmLEr+0eWI/se3O8U
aGH/ZjXd/Ii3bCltjbmBxHzsXRiAJdWaZzPnVwjJ8ZdpPOwuUPAXINjDQv3yGAatCVymhX5GibVd
LPdl+nOaLYsx43Zh3g8sCk3bEfQayYLJKObFvXJvH8/xPd2t4wzDW7320rKdsNVypAepLWHh5TqF
I/4aaptXTBWipw1pcbx2Qs5pvPeCdeZJ3oN0m5dSg9Fq3bVNXlJFtge762wkYMyPQwpvN2c2HDYr
P825OnN9oHQCEzlGJ60il+Rq23h4c7HUYp5IHS7v5xOstTyUyXGjpbUnayiV6FTtMy8bHeNibpjn
u6i/m0ehRP9xKzmlZ7hWzgUaDTVENehRik95R/9tKV95E0M5VfRU0VH5nK1CijK95kNMGo8yvcBO
FBWBTzut4kzEBw5m3YijUqfTyYuPaLBa2N/r8jG/Mz5c1PdHtFpv1wulkUbjE+i1bWL8CwOjXU6s
0nvorX7eenH2oWfPbFqC0IpomMYw7Q1MdsyPpwACxFQ9Bbm0MCdmvJW7l+eLrzipdNZjCtN/NZzI
kwX/h6J6PNv9ysi+G5Mr7wOvR0majjnUwGPfTSCtlGotm1Xz/uohNHd20W9ry2uj/RdNkwqNgTEb
FhPlBAxBfcEgi5Q71atau77CSYrpAZGZADTatcJcm36gSSB00ZVPOi19uulLRbgjYDFlaIM6EOz2
s0t/JJi8qYi9HhRgqAbElbF7zO/JqbA5Bl5ydhBlOGrfyXT1TeTPb8RgmB3E4zg13wvodBGBAE9i
/JZq9TCk9Ka8xS2XF1AtpIHZzA1JK5XBby9HTka1L2+QZUwqFYbYfPVoKAZTo9ekhni6+cGQQgK3
LtQ1MCGrsN/1pK/iQ1oHHzBi2+WMUGSalacDJd0KUigygrMmRidKKbUEtGnt+bw3Terkw/dJsR6G
ybIvlcvHlkUOv6un6i2+Fc4SROVh0dU/ZQ2FICTkN78KWaNyQEjPRQMQ/bHSG8HSetRyrrDnvr1W
yhXxLkS0gY28MWRPJdICFl+eWTCjMGKk7kZgRzDApPPqSdFIsi74JhXAXxaIMHNCNEa3anHu83zq
bHu81WO05mbxyaRW9aM1Cw9bLcHNg6OeGmW4lqMXc0ZWJxZao/ryYIw6JrsgWUJ5mbs4RiVap0Qt
Bwc6GYVRpjzs6X3/H5Cjlo0w+RACf7NGoJC035oqj9VIPOb6oxD3YlC8w7pJiy+Dq5dSZ5YJ8tt1
q1BALbWN0LXkFEvjMoxiRiR9nU+W9HEH9O5/d9hANg8khVx6TlzzLRydpAMvGAIY3kjSG0lFs3l4
L5vT+U05gPPrPPXgaQ6QHE6sx4QwBSW1LQdI+fqX+Or8jKjATk8S+wrGNOx5T61T1bye5+GwRsvZ
srF85eloFc6lnuDn3PVJlIJMzLGyWweS6m1bGRtJGfNsAOOlqD4VY/fcVhFv5P4JBlHFvvyIrl8U
/HwJl0Rs2RR51NHOqiMVDX791sIdbAtXUBYeYA8e5u/ZWtzfN0oHmCYi1lLS5vp+HYiW53BZPRx5
YJ/r0iCl35GZquAIyBED/9tvGtZKZimJcnXMnqtpmnwwclaIIA8Hk6aR69MV8h5dPOWI3Wm2fKvb
FpzKE1LyqjejtlcW/HnFsACAPY6WsY6757/bW9MxIRVEf/3skGP8QS0ESps5yP7JAgRQBJutzEP3
O8ZwRhwp8s9KUxvVGFsI6xWBD8j6BZDhZfzNeEKrIybL8sVYSJ9olUpw0dkQFhvtp+MO77uW9V10
9IRX2Ob/r1jsMjCCvGTZZj/Kidqev5w3dml1YJggUmKj0gWlIqdHDuR3VnCUSoxX5soqjR6sBM8t
EcyakjtsSrkjV8Bl1lNrxcSez5iTaiHT+MHp0jtmZ0ZKt4rMEsUTi6QdVAUnlWZXck2A+GMGDLyl
iXGDALq3tj1yZK3j0vehHiic6dW6AE3Dgs1J5IHdIP2aMQblRj70qFZDicfpR7uyi3OGbBqmmMTH
KOlr3xT89aq4S5p5y0OuL/iF3q9zU60AfeuhpwnsC7gjQVixGc7iCyL29vZcXyZ9s9QytTub+vYm
OCDIFvVGDB2UnJYGThiLzBMPkqUJboBIEFO0yayIBEtOhRGoRgJ/znXlEj1eb/dtLverbyS5ZWa6
p6VkinBaqSPuNjtqskSz8NCYeZGTs+BXP3t0vf/0wcavoGO3RbWxOJtbuXOdNA/b9Ruj3QeNrG26
0T8lzikTKOYkod5qRFv64VlIjC9mhKi4alF4LhHKZpqA16G29JGrE3Id2cdN6CCig07k8sOQqbTm
CchWh0ousZJZmjQG732cytgxk0PD3JlPBY/NUd68Y/10C8l1GCVFCMDI549Gp8JvOkONMzyfgq52
H9slLvwNg3y5Kqdm268i547LbHGOObpPqV3ecbkI2UxjjgJQWwHsEJ500SPiplf0OXKN/6rcmRGz
a4hohBlULebapg6S8qHQBUv0gbXJVepO2a3tdryivLgFoIX1eNjIR7VzuQ5OXgB75B3zYwc3dWY8
somrcBwJX8WRDHHU7Q6OQGbAaAs+D4vjLp5HhOUKkUvVNXja1YAVLFayD45IIiz2TwBUGdaGtqmR
/GrVq6uV3PjWZ8uPicNhdkZeEgsysypHPfIyowDC8JDveVnMWJLn4BkgHv34Mn9QOLB+xYBDtBxx
NKdzG+0nzfl1ve9WxOnpy+ULoly6Kq/s01PKT2ZPVK+Nn+zLGcFLmo+dRGOCdZt62e/E25FA9ocj
ee9XEjDgqpF/NhhBdiOQUTrpDNt0b2HkHw8TFtXVCsovzZTV6kw/vneemdICiGsxf4hx0wpx7bNW
76WdikKUoBv71ehjkIo5H6a0J7QJDqea4UmjbHP1ecrQWEEClbdVo8iynJ9la6cQfTLxPMqRrLTi
JM/ZYnlYF9KH+BEf0TtFwDYd5tW1YF6ESCYPGsFR68lqQjdL3F/+1SZNkX3YYAwGe71akPPehYsk
onWnyVAemlQoA9DZSZLRP7j2/qYnWy4Td36AAij+yhGynzlkvJY5pDW3HljduvSh6zm7rl0jpXY8
hhVLXwO1wR86RH7R3u8BUMHIZqXQW0kEmdcg+ZFfaIW918nPOdbUb6qvqoJu+EYsnINc2U7xZe2k
wFXTYrgOeN+YQDUJxFJM+8sDJNcz6FLy0KpN1Eqz1njJS7D7e7z6F6hVv/NKC8pxpfEH2YbZIIzW
OZFX4PQM5nEQlhtPb0RGg9KWkYun+FgcyvGK3IPGXVDzQH2hA2aRgNzCNX/+Q9A0lEvt/HEbEY23
yUmTTPe7pIDQ9QGabQIfJZwwRohEMXw63v9hO+m4ljP48Mp4yV4FkyXeTl3dh7yQKATM3hwX/CbA
hU8+V/89yMTvJEIfD8JEmQD7byD+Igt3LBWlfnj4ycJBZrPMc8Czjj9aI9pgNWEfQmp+1aBJhDlL
GBBKDVY345UyR2CGmeZwehKZ7a6vt2a0UDbWoxJvceHXAYsv8Kfoy9E6yWudWE5SHNGwqRSIqQzw
DHSL52U/S6NU+GfecRfpOzXDBg8U290PqDkIGCay0kot4PXjBvrjZIJ1czVb0+NNdPJw2Y1nfDFp
Tit/BVVXD857xQvDLc7+K231aPpHIt0vYuuBIwCgspoQ5976s+9ewCGLikSewOVhTxDGAF8v04oP
Qdf6ttZVaOB3Z7xUJs1wneO1P3mARUz0rqN1y9iVfAppuginPAGyugDZUn9G9OMyqMQ62SzlrCm6
wny10UnfPwgJM+esnjoRTsxrPsIOUGgnV920lOybYtD2XDaCvxrKmBRZhdcV0XR/mxAU6wQCQFXi
Ts+ICWBY7kxBIh4J99ZwlVbwaO/ASOVH2wndWdeii/qh98nvsmpANM2470Kv0zOlyJuh17kPTEJd
Aq24NDl2rJSYmPGTcXISXSSgeJgrJWyyOZpQzf/REB2RNEvbRopA92kW9tml8UXANqNZ+CuW6ByV
HT2hZ/tTdJiZYCKVakoyO+lDpI2uFfFLfaeL9HZNFDcBe+XqpEzNChOA0MpY2zI9pIlUudxUJ3/v
sxxfVc/AwRF8Fp+Y+UuC4klbP+ImUWo48D3U1lhQcaUBWqmwSxcIRT2ncLTbJcvyZRKrU1Ir1QK4
rrgSAIWhhjX+VlMe5FMVXvXQmCrQgrify+EaQFGyzALhZ0LNITYLuUiDAAVyWXJToCwIJDZ3Sn08
3ySlAK24jtIKnssdjDRmCa22aomNEPeH6bTK2LmiAPpB2d47uzp273D6/KHWQIc0UcxHYVkogpcu
yMtH+1C8MuT87WX++yjwfgJamvJ347PdsvLCRPu02zSt/Jc6wR4gQ1/ycijml0cYWKPY8853pIKw
mTGlTI/Fmqo2trj3DCPed7Ymy/ht0ZVspppvr3a4Ot4lhj6LxqRxlBky1Z1ub/etmud6egaHKgd1
gA8Nw5ENrsfJw0S+tr+uj0E2lzfFRZV3soKJc52VW9auIkDtvaF6hdd2RjLDsTwlNlTjfzwnameN
HQISCkuwS6s3qptXBMyAGuib0mPncQhR1z6slMNOmPp1ecOQK+i8MpfmDFnxd63bPIyXVqp3H/ft
PBoLlG7WIF9hkZhJD/unjdXH8ebjZGoyekn8qUSb0B+/o6DuYqmXvaKoeG3/21G7l5M9PfyP4MnM
fNw3i8IcFnnMmFm+/D/nWf8x6O0MC/oQbtpHLW21va+Gcmqf1KgYGOLcL46Vu5XHqRLA5Wa74g1G
C+gmDfFh6eYy9FN8iavNK/tDvSqMvyGUs2Ne50q/gd0MMe958fuF1jCh6TMlIJLPha/HLbecI8gH
xNm+eeGI+e/uB0+DLuBz3CqkLteD/lNi4TP14gEDRnkXwvCZRNV4BVXUFYCbJG0dl8u9xtFNX5s0
Odtqo5+aQjPVcQ5P6NkEQAD9NjoYooZdOnSAz2QAbnsiAULUUWa6pZn98MssJUiFJkacw42PkWav
iSkSpzeHYMOZFIgW35iNkBlWHvUtPjPu6nXixYJx02rX1rAJy8Ere/2NmXt8II2TjxsKKtOwF6if
yeb7XoF/6RZTUZqH7xv/aNDt/PqutBd2h2VD+ZfUUmiDYH9kXV5f6dvNJgTYhPnKkNOn4SNGE4/m
XYrAVZFIP+9vFAT1O7Ef1K72vA1KnIglgOr7znWbqigHOrX+0IJQWJR59OyOG16yndbH4oCjn4l7
0OZow8M/c5GAfDDk3Pi8SD7Lf+eaDLJmjbgotgAG0twtaCa4/W58B3hrqRRw65hr780jMdP1eTym
xPbc3S1616ahw0/g/F0lIYb8P6520cspQS0LnpDlZfNrLUUXLy9TnsCqwqb2Gh2+rBMU+Le0tFxf
bfaQiFHyOKWZpdROi/vNSne9rjhI153X/NiCk40vLRWCKmWV/Js+P53NnDWFxfzefvgx9VW3G/82
SFu5EPN/hF+XNFPfdkf4v7KXExwdiGkS3FyeRpveL/bdvcjPxH0QkPuEJhP0XrT40tH4oI5uo1Nu
StMlzYSwX0KHs1UP9suuvh1/B3pfo8DRFGoQqUhUWjBecB+I8sqPrE6k3MVzNOJXl/5+ZwOgVt6f
izJlRPW60A4GcJ0HKAw2wbRxBqwCFdUBxR1+/XAaswupRp3UYWWJHkf+3aHp7IzqPiX0taRCqVsj
4GuNaSXEYFv5OB7uI6t23nFFpzGzke30UZ7FANpLRYLnAGwnObtTcuNjkAAPgRq11ggSbRsTX77f
eaxwzZXGtrYKmkpvC5cSCvaYeXXkCsNU1FdiDGsxwPPTFs3PXUcYqLrqaiDEonMLORLu1Kbrsafr
cdanDQuIISfwwI3E87HVRIS4vtAs2yOhcJSc7mToeD84PhrVBin3w99GIXapwDj97iX2y7MFffjF
WZtQPztl3yV8jDBlaMrZ2BR2sP18ur6w4WTSXaEFw+F/dd/+4q+JbOhHUqvTu90MQqALw2nIksoK
Hj9ooD4p8wXtAPKtmKipxCeZBKYLX6GlSzzPvwENxodP3cntgAU6uXKvSymYqWZ2VR8MbL52dPBH
QeU+v7iSQ6M8cTY85jeo14CupNZZHfnWbCvTv3D8gFqyh9H9t1HQOcRtnYB5pKC/KMGsGvqlLooz
JTVULPwGRakkL594keTJklu7E35gm5R5s/WeiUtTaYoK/NqGE8b5LTuikGYEvG6OABfjuj4l96AF
u6RsFrYHOrgz+f+IeGgFid/SHt0nNMdutlPSdaGAXVtSbYefs79EIbOMRfsvMbBxWc5QtHXaCsCA
Kzwkn5Jw+0bXGzAHyE+iRS3RaaZYts2IfWKU8TJYTAnDnrp7YnULyxSCfyaeAkX7WMNhoa7gEoVR
6lXi7JcOEBqnH15qTo9nMNVez188iq9dZEKnognFfaUXIvG5aRMDLGYL61R3Ji6tRSt4OxsQtPrE
K0D6KCxxHZ4QqwU9/Hz2L6oHVy4mZDge1YeDYOyKLCMNcMnlZhF8BXEG7iUeGJfbhg/QsezGYGSd
I3Xht3eJpvj5L+HxmfxHCQZynjYeniE/VR39RLquZ0MKLDlu1fl0ah7FlZACyEDIWJ6emf0tznKD
sz1O9ETqJIFoAWNvIh/C/XD9CBWh99yw1qQZdCD6M9VbP8Xi4bFr+BuPJKC3YlrKg0K4HIC8c35H
iSa4vDsqT0n+fpIz3dM1p8uWO7w50rTC4oASlXRfIGTYqOgRzY0/5zBC+I3Kbfm0BM92crcBG5DL
Xs+etMtd2buaaffJPUIVMM36IkSSMsrpBor4ttexMVXvsgPLw2ijbGwXPHtQO398Mnmp2ogVaLhZ
FC62FPDL/vXkRkKtpyjkfRsasoSpaXcgHhKsd8Q329rTShxaxNEk0Ex+EFcaxFK2IP7ZH+h3jaEJ
rsVdGRRIpSXnXAg7ammJM8ozfrYgQi5oKMKI3ez84+aH37ITinJmLKBDKVSx4/guKFCUKNhUxTc3
eM2SIWZTPvNU4pH+QXRKXqelbisrIdjzGUyqSl4tH3Wsnes83nL0G+3hFOhKGyXAiiiEvpHE/hPu
CfKamqFvwhNa+SJd/7qp4Ax+Yu2vR7+ts6jZjjC0HRkn2M9nJaRLipLkmsD5SQV6dRGCHSxf/GDa
DH+7MJIfq6exdy82zhzf6vXWhE7UlIFWv0ea6jO9uv7AIjXXqjE6mUTFBfLVEcUE3X4T7i7atbNi
yyrHpJaixkkKxpP+06vVNawdcK7OCh4Tl5gRv6QzE4gLUiY+D3d1k/1KDcPjP8WOs1h3LOnDJXhE
7PwBYh4YiHZafZ3WC0keImptt34jW7d/5Rqg+Ou1nYmDlePZEGczmAuFAG0SQN/EpzRp7wR+XaDL
VciQS45YqMBaDSrwqK4n2Q8v+KRRk1iC8ChNJd2k3ThzoPdnIBGHeEsVBZKd5lLVgSyHktYoIDhT
4SSh22RSGDGmjYHHl3n1rrfD+ZMr+r7ssnvn8o/tOUUhfIUhddz4yyfpEBtnVotRQ0DcXs2j8No2
Pua+RGa4HadVrY8OyKnh+YTy0ABpNtshvPcJeyL5N3120bui/dEEtmiyuuuagj/8rgN8fhoEqk+t
QXoY3jPjLrc79Uxy4oQBy8JQGukKCk7iDe5Uqg/EbFXFhuYLxO/2EfLAFYn/eqavSVC0XKc39Y4U
iKwdndiNGLEuijNB67o3paMMg0tvcFK8z1tYM9lF4NVN3RZbctIFsU629286CRy7NBqwb94CwDe3
UZl+nH7UswHoGzlNaa/032+KKwPc4uTO5APBNAncqUxi5V6lc+L/36aniUlvcPHdja5OcdhnjXKH
u7xB7w+N0HNSR/z3bnPl+u00DEiAI9gSsgJhf2A+O/8NNW9PZsYIsfye/M6/JEhj9ErYQICrf9Ww
c8wK1qMXzl6J/4FqzNZYV+YUS0tOQIeRexxZfYxpWy/xHNkmd+6PkP2uChH8nF1Qt4RY5LZVwA2Y
16sOdCiqywvk9SvtVULxtO+85OR/aHzr2Vol2RUfbTKqWXA1I1zBq1zu/fcekqRDtSIEZnUP7Ukh
iP7T6u1xYW0UnRQ3iQC76ko2VRwfXYIFw3WjZNptHr9p8L/eY+wS7amhoBUwQGmqmTAVxaa0XfdE
4AvZ+MC4xwZPGnXImN8Q6agBYF0DBpzQnwG+vxazybRKUbEkCyZovUnrJpX3oIzLUCuyiv8KDHPV
Br4EOfsG/UNfSCoxcSVn61NvXuq84BKY8WYKfkZKBovKZm/nEnAU5uTUZ7jlbusDQ3Sxk/Sz24Uc
7ejup62/1g97JNLSp3cuTbsMmKs5Q+R/uqF70mhgFNYMlw1TFZ6TjozbYa1JX1CbaxRtboFyal23
kwb0bxSrUB+JHLveIrr7yd7mHQBF8vf6+nDP51fKDbjwyq7flwMqTdjSBFPJgLtykU5hWmxs4JFA
8DEKMBSYaSkSkfmZDUEmkP5HAvrGuKhizjNnmpaboCfFXcRrpa7hg0m6bEkIMg65VStGRznp75LK
8YiL6hFaMBSF46hKKSA0RSkcY2s98apNun6XwLc4l4smP9/BK7+VvnaibSEaksihVEITURp6Q9Mr
7RWmmI8OPZaPMTS5/VZ0XNBSFmd2KftPsm/4mI5lT+1UPfUrzkjixsBl1CBxBk0+2kxxdhd2VGMO
Q/A/3kM4tbY/wPApWQ+XLfxCtrLIOg1fQsgwdZ/gQJQ4KwLU3wrdRH6uyr39cP3i2XbS7G3V8cj9
DO0i78XFoKvnfNZP2DOUYWW4605bgIk2q1YbRbYLx3r2Uf3hmue4xY/0PTZup8mtyz1IMyBKhkYt
9hkRoqLMNWilRox2jLIlzgWtdqMMHPwkVw2DCAa6RG7R6Q4fTfJm27uq2s3PtcPbbADQn/452nij
fICWChyc95j9g5kXZGNhC7V4ToMBn2+uoIvrhFamNSEQlvIFQIPW2FZ9HMkVxnJDhj0Amo0SfWAr
4ACwUtUaQe+ZpLDEXGHiWlD51psJcuV8GVPVrjy5r3t4fqR0gap3z6VyzkMT0XrIYFNBeGHnSVjU
0pZLKYJiTMkZkttvQoMQokxPa3+tVwR+km68Z1dWgkY48B09SwonhR4gDDeKn8UyLleTBQiWZUKZ
WPyCqe0cIY1TF/oBmnqdhdhVm0lqXbXUIti5cexxmDfJCU1LZTqcaxXW1IS0+qUYvYH1zX/fcyev
BHrA+YyE6lpnITz93gQC0glNFOqFtUSahPWYq1E5pgCf8wPRHhr3HuMTdUKpnw4fO7b+eaPITdNO
leJvu+v8W/+2tgtdAQuyFinxZ76PZzI0IvIxlssv20Y9eU0SzuoLPh/GzmzfZ8sMvGGyckbJZsMu
G0sKuEef5WWQp1x5tWkiQFRgmZazUAGzEEtDguWz1ftdCAl0O/So/BstYDGtluNJr9nP2TraOrcJ
6a7PI2yKv2RTHzrEf0Kdy3jR8xlIEVdnxJGubnCZGuCcm47boJsQDKnax1+OJFOQCCE5tFfSlzyC
uZV7Q4zMG7vnOyfDYD5uhXFuhSj/NQD5J/nxi+8NxthNponta6HswHVIS4rrJPQAQNVJ8SezMwIa
8KbnZm34vxFE9WTluNsdgKePnDAt6B6DBjS34OGO3+pdf6gqYcFZ4qPhmzWT+jBghCXmyDAhPVtk
+GMMZFHLX0uFOWRDjZXYveXVMdbCbyS5Pp36ciGQCKUze8bcIgCzcBkneJ+ynahgqE6lDhb/5cPM
2lSFECxy7KdaDFYPk6b8q/0+Puuzqa3t96NAMmyLxVFRrvHoAMxX0HDLdyRumfwN/TA+hzaVk7AI
wgaQynP2/NlZxLuVH+7cOBqgbUd5x/z0iRCCnLZTXL+9EHvA4xF4TVSu9wSfXy/10/cjQ08uEhOG
ZJBOhObqN9vXLvcycoqLKIQDeDx6+MX4VfOczl3ZmPeWBAgRSMa0eNP5/KNHp6K7pjA/Vhk3y7jh
FwbYS0uwCnWZoMlMq1kzqmnRYA49ysbdv+S+wNEW9n5KAbCxzHx1fU1R9QrqjktDi1KTnlQadAmE
UHaPTWDA4lteXFJdJIOqlTj8PYcZQsJYn1vjArwKZM8YTqTJckxlDSgwH/PNFWA3PAYZRHDEaoUt
vfCWmjx+U76jFhlwSViy9hwDEY1HL59mhYYMpv0ai/BmVSgUHUGWVlPUtVN8DHSciVT2+QBssPHK
cSHxn57jhKc20hAE0fo7dgXyy/p2UpADJi+P95EKZH31F83gAGvuOrkPWbB6QYja5RxgUxOA0dDH
zkMnNVnxx6n5oCJLpWMTRgVX/kgpSafEV7DBZJHOS5aILRy9NPCEz9GTBMJGDy6ekiZ4FUqxWBwo
I1dZ5Nv/9hc/Acmc8UaDm8g57A3VQ5KobDuWT2SDZTrR0MPmnF6KsTzg9ulTuDR9Fc8EFKXliRL0
1+IXKsIiK5nX58Oep7JqL29vLmDaBMM8eqkT8qitbruTIZ9rGM1eYEv/W5puGi6pke9Dx3BjWyGi
YQyREzEI1X9Ev7iF0jxtncU1CUP2NkNdXrQksBm7dSwUv6QJDte2Tove909rzG5rJvCnOEM9Lxk2
uqOJTofV721qGoWGabfgXG2q7YTmZyvdI9ZS8BRnZfPRvjfAGIWd+hFuahGjV9vNjhtS59HdWx/2
w5J7spCI6/ZgGVVwzOuRN4TMEtmRuXhKIJWX4W9N2mmFD0HfMyvhdLXwDmR5XUlsdWYkZKt9eY/V
auVYcho6Okq+CoLsxsXiKIjJoXYizgwG3Zy1rt9hz94zqodCoMWNvXvBLo8lKXAjZubzutPnzx8i
tJ3FaKhthFe9JiBHfyMgfJu+DyXmePdSs5HF3LwSId7PxcGQmx7hdUlMDlz8FpD2Cl/Jiyjie6Bv
cpciUesFAC95Dq7oe+lq09X154kgwyRjLQPsc90IzDl5dmowN2Sir0VG6bHdw41uobXEe0t2DW5j
iaY8moKA1pChGmTt26d8psxi0OedMGNifQ5MCgiEgjW1grP1jdNsaYdbnXzbNRXeG02thyw3IqeN
Xf3LvYKfOO3J0CN2llnKNtGsWyhXrc5xlKRQMlaSIU7Z9hOp8vYhJRrtRZXIDulCMnz0EsezJTZj
j8Lnm8h/yT92muZNHGmjOk7hIhXClBgKZ0CqNPEGnA7vfkw1GV5FDwpZBe3p1Nq1+YU9JEUOxyoR
xNLbABxzyNGljom1A5y5O5ikJUzTOZEdUG9g5zJ7XwF4xGtcMoYtrFQTKbo5zkNyyblZrimtxLWT
BcM1q0+PVZ+JUZoKsvS2W4DslE2nucGGGLbBpuFIF2/kpU/YHtD9nINOF//O8Pwt0CRTiwr2LBPo
UIypck2c36nSbza2ReH8AeIGvF0Oq5S/mXxkQZ4lZzTSRFkVH3bT8V5pTRKsvSWV1Im5n5SGuEA9
o75SFiTXy4TQRcwWPIp+PAYVjCWJ+UKDm5dwNtmAcZZBXSHI2UY0WbPiYYAvzOYFq9d8uYKRE3lQ
MKMx9sWjhIrpY//HtXqnZNxO+TNUHZBOhjWXY+tG+UBp3CJZPRM4zMBemyRCRqyoaIZakXy0K6zZ
hGWtAKbPG5mvTmZwuY2m2mipwCXRAlEXrQ5XkNlPwCjpLQhCY55TtkTC0bXiq7zZYZrY/bOekYLF
gE48KQoYJA8E4vnyevW8/9uCf80nCbX1A4dYAEViMP8+GYh5IhVkIxKzSA2ovxEfT1qj8bM9wpBG
W6YII4v4es6oxnY1Pd8fECl51I+5aCKEUbrNChbS2mB0As5rootYdoA6mTFq5X2+wpmOJTqun9bS
ouQ55r6F+9dXvm5GVn+/o8BujV+/ha4a1OLO6N3XhBpDTKrCbd8J5uSUQwaZNyvkk1blwUoxNHdE
Jf9DKj6OufYVo7gX+SnTvoHzgIMocBlQ/c9vvn88pg5UB8PS2Nvj2Psb+5rwN7/uMW0Cfjomxyrs
B4UHTS8lyo/xF8FYzvSmlWEVhzkdclioYILHLGYfYhSG/4JTAx+InZTHD2xztuPX1INzO2yUCMLu
WIT6HCVazbGiFCWf0KhsYwDwmcButz0v3cwPD3Y8oqz5++2+4+BA7G6apO+iAri5ws0QniIiYxGN
ehPBqEuhrA2MbhN/vNT5EsL3qBJVeIeaBaWV/3vRHOIVVdknZBN4eNw4jl/xZAxOYIhIOy50ZBy3
9cHK+Kapc1ExNI+tu+rwEuqTMT828GmLBnKYPQ5L4kex1SKYM+0tIbq2iRxTKE1/g8/I544BJeCL
IrYCW8Kj3SN/HDrG2fnLTNNXmzKw4vU8/3umz9KkuO0UuqUtJX1FS+hwsHLe/1d0Yng/J7R1C9JN
G1oaemTbxKODcATsY9eJn5xTrtunuuJSLTIBlvGWcN5dUpor3GTmnen37IrXTKT2Gsea7tGSOZV8
iUOG3HWY7Y6fsZhWHJQks9A91Yz48fxK9u1aRvZ6np6/mtfiZHmwJMktb+NFBDPGNbEnw9zZMdgQ
vl+84wHgb1NRXJUU/uasQKF6MXQsmvfiRsp5DDI5x9IxjThSC9hg3kog0E0lWvJvawleuQQjP57H
Hsh8RknOcHSfqnu26odAq36QqWxiYb8rhj/Ft56gWkCHNjCUHBAFUEYNinzVtsD8Ju9VLOMDq4LN
s2FVjZDBhSHLmjYYXkjBRuLNuuOJBYzJWSrgKvmMmpyGBnaxaRucMbAicwfX/9eq6dqWunpPXdO+
xi1QUUbeqO3Niq3V8cikdojEBPXNsmcArrADDIE4A0X95kYvV3TN1MJ8ferVZ/dsx3pOoFhpTdSw
m6E4Jc736k4TpsRKmHO9UZis354Zdo++F45PvwM7XWRs+l2KrUX9kEEzA8Vl7iMaI7QTmIQpwXDr
pVdrI46Hy2sU7FLmPinQYWdWHIsauIa3IWB7WF+QPbSnhWk98QRpb3uKBKYthhDY0ai2YMeoO/9w
zYxNQb6wZ1XZSeA7AtMyheEUQlLLcy9/p84mPvivKhkKclF8GycQqK5Db4WzkFa83j21uzXhMT77
sryXwE9gdyUHzCafnkcEVV5DT9YrftBaEyzzvFX7M6jOD/c35/4HiSeEkr8jBJJKJIEEAarr66sC
6V8EnFvZxECymbDpl9LQ5xTyUGZg+g4ABvoYkX7QukRsasKAkhiEqH0XUcY3EEgaswLY1c9WiPYD
rjvCuHCCAFbmercPgablVzDfb0dYKGnedP36x1n+l12d3lHbTj+BlnjhbhiTm3Gd9efuKQrseLcq
2oZisQqIhkRqOtNFlaLbZSrsMO2tuVVuq/eieYOr+oQWY+6o9I9/iU2EP/KwiBIGYOmHBl8yiSoK
owCysjauGdROs2jbTCILkYn/91tvWfyGUIPNwSJGQt7OJ92OzARZ6zW7sYm5dBT4Pmey4M0GLx36
DoWyyhr7bf3ZXNQ5QuDfTS/8+oulksYIHH3IYC7sgXxjqoEEvOAJzj7Bl1j4dyRP+Ew3UPa6P2GL
nDSlUuE9ZcB2wsPI1a8YwEkMdN40jN0KJ3lbzVV/+5m/qHa75bWoyxbepFSaRR9yI3XbL/BSIjiK
WXB2ER6vfjd3jq9xjc22SpEGyC8Q/VOCHpX/w0/64IiZZ3Yxh+NlFtgig/5mlP1SikTUlJZXOM0t
ogE0nbW5ZtJ9tkizSe1QMyS5yJ5DB4ErAE2aBpILCfLJBYpKZzqQPqBcAXZTcFqPfX72kLbt5Sm3
VyuxGKzO4Ez/Z9vQKObTmry55P2AsKz0I7Pgso/dPeM+EjD9y22ifhI0RujHY3HHKnOGOkaU6J6I
wZf1qf4lOg756ZLKbvSeXXTHM/O2nsAQYmylnCRRP7dZB4EXyjvEluncUMbO1u0cbynT04RMokRF
eLEam1HkcEwxRPbK04l/eN69SEExx8If+/tJ0zYtyrBRlzbyzWqT/XmMhvZtmE5F+E/9i7qQDixL
qbFnlbe71EJRekQCYRTMMGGSoOLNJ/V6xyYqaqC+0zF0owQFNTSyFfsyO6MMlQ5XC1qkPbL87lVh
wT4vPIX8wfnt4OvzG+yfp/atwbk+gjKo0bz/XQPZeEiqAEm6MH3M6Kcpd9O1ZpLluOse70hjfziC
xubo0JNsktcQhw/45llwEQvvbozp2oLpUJARhxHG+Ysdm75TIduYZuoDEtqKy2MiGdX0UwhIJTzq
p93syVCZ+HCuIajswYPnEgKwBIgzZ/JCHuRJiJtfu/DSRd/Wf23jtq4Y/AR+CTYgZlH8u7sLEwu2
JI5+NSeWibYxbyo8cxjc6lJiZ+Celxuwv3KrUI2Rz99t9sCABcdPNX9iSVAEmbzw/tgAL9qoRJN6
6r04iSXqIJ+XuD0yY99Wo1eRP3ODwrw0b9Z/Pk69UPOjs4jg5e/lCdbFurWLoVosFiVM7TrOfhD8
Lc+diRbhdbjaGB4oLVS5mXozfHnPjqzbnNcZJofIFrGdCMzMruN4kflJt8MUgR3uu45Pun6xKVqg
NBN6watq6ZTk1ZGDF1GzTfAmCdOUfLjDvN6cpI2I2AIt4TDLsrwCih0fsReTqgPxeQBsDn7wc72W
BFK83+XvQGaQ5slW09dogqTfeLT/ICpq2vAkQoi+qvs8pPM5UjSRIPpHCPklIgiKx/5Pp60GrAhk
X4u0MCCaWtVoDYCO35lskz1vxU9+2Z519FQOGHkCv2tZTZLfuTtAzooboqZYuswcBXeGKV206aIO
A4ihyWVrUz9h1ME2p76ixx89xaJz1Yr6wTJOggLvDFS1BxF236/vd7zmJK802p+B4IbvXLgY4B8P
bCkOg2EaBlLqgQmXheBhzg7WCWzpQrUwdBBOUGqreH1ZmFUOmHlQnUx30SzK4BUTNdwAEB7chp6Y
oFFzIs+O1+8EpP9VC8O05DNcXiFsVDGuK3z2IAFEKNwPWM/O37FjU2Zy8aYxHgK/4On9YBgz7tYJ
yQUroawp+IenQcIE5K6RMENmYeC6qg3xTTspKUvmcoz19ukdk3rcO1gu83Yk6iBO+QErD7U5EQjI
maf2jLZMCjhUvEh8GrHi9+1LbcZz4Hsow4rhxGcDeW6ES+K54b+Xz17wEjxzGgPxTbAAzVHsX9iM
Cq9ZJ9wUhMCKgrC4FS+kd6uSBfogdZfsgPmRNxZs60cobRXJc23FUQUL+v3/stKMpTSR9c1MWthh
zVeUrwp/lV4K2kIVeVk8HZE9nNzDxs2TTk/mMu2hG9P99N0FTfjN3vPabDUusNPpFOTodqM4piOK
yAvtVJVfCCB6w234QQSdz5s5vVC6jpleuhCfc9b+kKzez1/lgOX1CefEdD5ut1ERMbGuUmzIo+sH
iZdFlnMnHhWGqEY4B6cpyWai9A9zPYUBiKXu+u8iGQBksjGI5jdgF3fGVNe0fDzYmFQY+exllbL/
F+1b1h7laIp3zinpckZAAxFTbyW4NcVakAKDRyfdxVwV/qK4EWYpTnflHnVn3xqMyXUosYYnWNSR
q5m5Y7zPXJYJx2RrchXbaNEvGlc2m4ToboWCVv5Qqslv/foYDMwO69HmtHkBN75LlZKvBGppZAVt
lG8iC/zAbadbf7HPAIk0fvuGIuTL1fET4EVP8FlX21Oqdv191MNydPSY39Cs3vl+AzntWqD3Y0mc
bI48B55fbQDFvajRAzEz7VWTkGMHO+2EIF8kWuFA02wJhd5Dvbc+jt3mWLbQoU8zVEFdgtTKr6Q+
fQYjtZHH6UKG0ILLs8aKPxflv+2HQaqr+pwo08yV1H4tYOCYXiLGD37wP/fRykYovbR6McUcdfZg
NOv+waPA/0pCxsO29PpOI86MSwGEbAYidQRO633mKB3Dso/eZmywgQmpzxjPCIe8aNLs3NA5Oey9
PfJ4wpumeedbkfKaGexsoT3OXSpP5BOUI8Fe5tYgxlLbTqxUsFjKUO31eF39khqUV8hMliPWdEak
v8IMAaKbcivKvlUMgVfMpsO2JVWUUfVjrMfwj+N9xl2EbbE1zo8fotqep5HEDKIFBNbgObow+QXV
t6CaL2dhbGWf90GZ5avvJkLw86CC1cCTISB0siIFf6TMURSfFkI8dcIupdwIggwKrylmoW2qbaCv
cSak01XyUneke8B9JzBhUC5GCsUvDOG4RpKY0Lvbg30NLPOL/24BpT74b2eSwR0L4JLlyddVykZQ
L8KdFY0s1ko7VWqxKInVPU7NtFTgqJN8kOKG5pNWnVIcd8cwFGao4gKnvQZft5cRmCuhowQIbrZr
tuH+32k88fstMW9m1q+0cRvQItakQY+j03KcqQgbb6j282Pp0pOUMKWeeTn+mPeOZ0HvvNtI6J8Y
981HUNR7JsQG9HIzvbSz2tPsP87FNLIZ0NftlyU1NNYE5fs5JBzXmvSYs43A1IZuUweDKAEdi2r5
9PktuYVxNnjksegnjfXDQkh0CR/2RvSU2aYfLYYs0sDvPDnJDH1Qkuh6RIvxUMJFaSnb1hprTgGC
ukyguuO3Y7f9kAU/KMImcEcbme71XZFcOnYeKNLGvEVoRjcC2es1d/AbEm3eZNPr9Or89nkBghA2
rf1MRXgBWFXwwOZG3aoq96qP2L7RZzYQ0hES4K1KSN887PMfFqZfHBLau++ycZiSBrQ+RQjVFGsU
LV3Tpsc6O/xXVecQQOWF7dqyNEYnBzx9W9EQ1486Moklm1sxznFPc2WBOGiGPn9GFjIwwk0KWWMJ
xSESe7CCyLct295z4XRh6YYYGiNb4Vw/jelwmiBZVsuIVBPozw1j6zWVh/lZe3UGvxNyoST04LYa
0SYXWiZcL0Z2TcblyaP364+mRcDSZYSDMtYo/dmWi1IVr4ps4wT+R569T64B16wOUpwzrGqNeCRs
HxrEEeehEsRGr1GNqPOKyBULeGglDqr/HOmH3+BKilBXf5xLr5wMNFB4eMAxy1Jo+diqpnN2Ydz9
JrYO4We7osW3xAUyRsEW3lXDS4Vc+xkU3DgYX/mbRQnL861TkSnF++7AVZD7RMvO8nSBHGqnKqGf
p3wPtP9stTTPtukCLX8FJyOQjY+z6CjBWPierAWuUM0AelUfE/s+DfA6jywDanN2OOZW6OjqJN74
dnG6fgqClbnnVTb+ctRy0vLLDfAyLSXTXrLMGuD3uk1fNTj7f9ELerJvgOas6ndh+JDjIqmPZu+y
Eb+vDTDiqe/ykt3cPIQICf4ogP5EhTXuplA+H5S/GnUkWSo/XswRw5zflASXAQuRj1Mt99fIoRJ+
By0KQ7ja0wffUzj9dFB21GAukQzLKezmdV3rhXkNclYRr8PuX1WZ+NXEGfVeCrgweibe30CqIBbY
wekfRMe58Kr0QCJcDTP7DdSW+qEXBYg6f3OmFJ8317GJhm0luQMsWDxpKIsfdim3lHDhZQuqJoqy
JUfp16YV7tE8nb3/rudhjlaxmOnqgZRo6bSa8l1c9BrrPjps5ium74cnrMBfYRBeySvJR2i1PQDf
MXZ6lXRhEe6qqU73Bx/BmflEaLKtztiEOjSqxslkg2DNldq7r5HmFhXIFYluRWJykTQOWA4b3t0e
q0M3bbcO/J/I0Xq8pyBS73d34HhWqf7IO680pHhV9mu+qrWk8oiM3scfyMVTwt7NLdJEAw+5Syrh
lLcixMFpy7q3JpTQ8Zb7wvQJZ2wOuqEafJfj2/tsf4rfAMu83vSRErSiKE45JvQ93Equ7n9QYyOV
QVHLzwp0FvMb8CTsJF5gwdS2IBZVnEXqBL+teozXXX4TdG3UocQwMwbBFfi48XXgcGX9k8js7+mR
vYfEtKM35+4hOg6xyS0Dw/BOTM1K66FiThpWWD7iK5x5UQTYO7Y79tAvfgMlr+/N4dhSzRroYEV0
ohPM7od3B+dOA2Ad0MMFYMzl86+zi2hLLOQpwSmKAAXHrwHytcltduYZp5sSzmJTc53bpLHg9EXG
ZoQQsd+oFOF28ITOZcgVyJPGgExRNNyMP89DERrD7nTcH95vFNTS0s4i5IiHJkLHZeK6yWEuCQS8
IOKiEf58Bhw6arm6J+K7HhEmml0sZ73I8Cu6BqNV/+lebBhMNksuIpEdD8lT8P59ePKZMp9O7r4i
G9t8Gtvyo5Pu3te6dV61AKJiDToFrfdNdgUi2ouHb5oX7dK82+9ln7fLR8aaW5VM3QpSPGCcUjaQ
2FG6uXT3rctGxXJG5rjBg/Z9saEYs+t281PMbUhG0hxUDei51B1qEjIxUjYt41ZpTjlsV9qBG0Ft
+UX4QjbQn/azySe8BBOTvWZ/OOF3dzX9KwukSUdQ2FN+YwHon2GYw2Vy3JPJTS4Gh0lRqvCBU+tp
2xdsHmsXD/Y/WsYX0nIEsxzwR9JNDhbVMqPuiXsaDIDfg7eyHD4NDcSFuEkQqDvclJMh8ghlVC52
k+FWP8sZMKIP7cQyE5d2Lfg9Ssgq+t2AR4+y5M5ZfUqD0QJRXetQK9G6LbQQFSQii+Lnn3MPn2rz
accWFyX22da9taeOb+11xfmvoqHBLQQGl7rYAlHZEINrKRBjoZloyPwQAS0LH+W0E1Bh9PGI8w0j
3V08qYfdWv+Ijg260TDTlplM7iXbI9rwrtOmusQN+YHSNQI8cd8bWZ0Q40ulrJEIXSxtPjzbeH7+
NhvxvrBt6ZcLaReD5+u7Fgyd9BwTtT93SI4cefEU6j8ymabQDRkTYA7bnfnDBCk17Dmea0Sc/vly
Uhzv3jymmYOhe9IKXn3keazDIlZgV8Tct3pniNNR0VfvSkRMtJ0gHcgwMB5ew2DLI++oMaRCs+nk
sMuiLh+WjLNCAXGBL5Fg1LK50ejIPHRmYgXfaIIxhlaCvYtp/THZffOo4RA4CHNO97zv88cgHalA
P+XYdD2uIFuhUCLU7h9R85MnboCkfo8bDFKpepFSnNqCp2LRMSiXoN6uznWbQOyM76ZH5RSJbnUV
Yy7vD2wkTuY7WoxXxsOO0tpp36KM69L2jF+pQmN97qo4eCUBxKzOPWE8iU6dI1401z3+V4HgzxRz
0EaslRkb2TSWyOXhETyHbd8phcskTRK9raRAF6SYwtgNPpiZI7TnhhXVOdx/QXvXpC6dUye9xAzl
VPEjJUV1lYx54mERNfkQ1HJcNJ3Ng1ChMzK0aqFv4LxD8GSnLvuDUg3wmgW0H6/FNdFjFYzv4YKH
xEQ8us+CabyMP1+6ce7p9fcS0tsKjEHdiO1LtbAaM2mlAbUR/fmUe7424JCjsxz6qJkVxuhAZCRp
2QrDY998/lRDNzJNWAeIBvZtFCLTeGkKo+7+ke8s9IzTjX57XA8xrrVK/yqSozTZd95b9f+SzZ2k
sJeiw/IOwVL05BJYTEEqDyMxAeM5izOBlnismEsxdLnO7T8pVrF585/aytxCd1C8JhL2nX3ORv9Z
Wpj87pTXSa0b0nhhA7gDwd9xl+OfM6t1wUiuHOV0RdOIwCHt/6zdr2YHKdBzQx58M62oZzIrTXN9
VdH2ttR3aeyccUBTyTa+8dMSZvT0ZZxRRx4B/cLeOJ8E50M9TgQ18QGzPO/MQQKIJM+YaAaIv+WH
hHxKLNEnWV1E1hT3/JKs0NJA/ApFugea+ojq4UG1ZMRlUePRex2boYfdzgg6wvligXwuTVNlhTpY
ZpvuDqx7kjiIKPkN6110N+fH2gYCXTftmyRoNaEXC7VEWq0t0385txxF4k9N+xq41Y369ezEl0z0
3Y3hC7H5Ou0GwaOuZ+nB0KFF67CIpmCqZnVM2MnPDak3wtXe6OOBHo4umjpkvCLK3DRq3TnwdYjF
1S6tMsrRgNdv7IHJAuEiS3WKNG2Aqjo2FfTSH1tanAAS/neFyHlGdDu2WQCdhXpoLh+8xDq76mOl
TuVBoRu9xe7W2PMoFEiOcEZRawXvTtdmvW7e7yQBzCB55tr+hqTVAnQxmhWM/8eBymlTAwzQv4DH
TpErKvJXT02sPtbyMLRCek0HMv0Qdv1Irm6HQh4rtH20Ub9f936RzjGQjZh/61nAR+L0VUPGzA/G
ua9EvzN+bXkxZKl0vfRjic7XxGS8ydyW+b4zhgB2snJIFvH+hWQbvJYQSS9xBAfwyYmHeqFGPnis
0Ugjw48UXZMtGSqkPeK0wayZUv2LcRvPtyCsUc6b1T8FVXe9d4h8edxrd/+hLFYQZSi8iuh0fmWW
N5MV/4CzkGbfsL53T3AQ5yvqlRHEit0RlCsn2kRa5X5Mt4MHn6PW9eB95EmB3rbwgf606SFCyGLW
sa1YtEExb6IJvBYfSfTD8j/7vFPJVh/A95cPtWd0tlZCo2GgmRks7w1OK4YQiwx7qwkkdcTekJqJ
8lu0/xeCzMAiu+OW8WcLPpJ6nxcIl0jmHTBIxx0UmyA+8HiOorUg/R9trWwqH8Gg/JBDrYlw8BVK
9pADStVRp/hSbik30mYOyGNuqMF73cwJa4o2uI9bOoaJnd4xQOMX14/0sIZb8fzMncVTS09eVKkI
/1Il9YkVI1AyjYd5122zD4U+6UrWrycMWwGA0SF6B/ZArX/4SyVFyXihCXP8FtBoFZAjBMnWwDcq
vO12kwTMjvWOjQNEUJZBYCdp1gOnkn9uJy9mSBINwXSIqNZqsSAsVZADK6kUxv8ZcRi+7mCE4X+e
FvJD9kh2FD6NSVN2oPLKUH7L/RB9zN69w8iEupkoLVisf0i79WC9UWG6fy3ic3eqcFGe/NaeMzr0
civ6HaIE8d+GBnV/Rt7DcHmah71bVxzaeMgRiM9uiu/2CsUp2B59ae/cq5rOFaCkW5B/hBbqR+KR
PzvOb8b194q/uwpG8OxV+VkyoKb7SMLSQCibAD3o46YlMqEMKsf3pjpIiGVq2XinIc+YlOFi0I+N
23dhnSqKTgWbYe8OAdDxgbLP/f7HkpjGV9zuut/YHzNK2bqUtjiqqa+LF4X8hv4O1e2YWmOo09Ew
kIP0fx/ek9/zc8UJ5+sW9eqn5goMrhtBIaMtNAXdP5uu8VZbYs796RB7NaxYV5bJG6HPoeJfbk9L
F4JA544lpWv4w+Wj5pN4LNtArR+i++psuhW3IqlDsbmcKg+lNH0kbPkvomK4/x3w2Xdtp61bx+me
ZkrRtp7jE74OBrNE4ex/njFvq6UO9yifXq1d8Saxtluln1xp9TZmo26ran5Ge56BjP6CF3serQk8
j9+sHlDXZhqU1M9gsFrkW3IfZtotZFd9UeWwhfzjQMsY+IL9pjUPo2PrdKZacF3jg42Iwckhaw3N
LxB525NYkkTqFQ1aBHDwIhhJ8exQwEDEwW+KY/56ANKNxF3lvbmui4HXAnug/5K+PrmEOZ5RQNXi
KbdIh6eNKd1jSJGhgulURDkTpAew+KFqvLx3XweQ1PlbaThAf1Za0AVWkM26RclzGVnWIkAWrtx8
sg7WUS3Kipi59jfw+iIw4Z5Z1v4++I6D76KfsyXZ9I6aNuIm9+eB09xIZj/0Jcg/nEyM0oD3N4R0
OG11ZJJS5Wq5ADFiYonhGkeCjJOOybwq7Bb29PNOncw8F+BAdlQyOHT6/DIBaM9dx1kj4jWErQUx
5FPHx5QQ8vgqrJzAmwsdTtFCF+kLZz0vxwYd2rCChfx6gD+p5Y+qp1YQjXEo/diazfu2jssV0C7w
NMWQtRt9BPOUHF4NX4XKbXTTl0OOYXlAEbAd9av5akcbOmBanvPmub2Igb0tL4WBecpGrKcjvj9a
p7q7iTJ2G6Um9dNYtrEwf9Pi/C1LnDkZPFa3SwAllbPQ0Ra5FAVMzYELQy6mfu5WkhDRyoQDczXX
G2Yz7SCwxQiUonzhbTDs9YPoNfwl8/e1xvRV5JidCM6rgGNavzYQ914g6Dz0WyEWUbLJxQ0uQX8U
jxaQeDWSGErwCUosP5BKRzK/OnrF8H7smcYhlVYCwwYumo7fSZ9ten3ngtuRofuid275VO7CfkIj
BCWklHUaw9/em+6ION55hXPbvHeg6vaxOZgYrLQ0z0PofGjM/FFV1ZXmBEUwOsXLiBbq10rw0H7l
Z4MMCeenPNMhoQIEcYdEDFf97wcWKKIficN/tTjFtE5JIvndrUDG7bNKGH+2XPiRRlM8x/L9p+ez
N7xtRtIwp/rW8y0ok4LArZSLLVm4Ly+DmSGsPWPX4qOKunZbl2OIoI9wnhvL47C3kHtE5j5a+CWn
3718yXdWFqmcKwrJHrUUs3bb2iqFNTCw5o3Un3YeJhOZpo0dVV4GsXic0DyFrjVGmxFOCNEkqYMj
kmzgYV7VgIEWKlSZysfFMPyPKe8eqLZvf7/pGleoh1GyNQEa2v8ZRHfebBfOZHqe/7Gubx/aUint
qp+GNA8LLfy26ZXhjcyN8TLN23mvHuhYSBt1RJYvhqP5+GcGl5pWFLMmZJBC47y05esYZVNZEpvp
iF5lX6exqCRUHgENWHOaltjafWZ1yji+DOAIvF55COH9N8TpVa3W0P3HgKg/oncF1iPi8bG3/r4G
rjnwz+exmIWRQuYcQryT6SEd1CnUYZCYQSDpK3XlI2jzObX9y2XlzhTvJa/wPJuO8q1wNlzGe70T
Vsxj5Sn+XdgzX7EHiG1eRVTT162770jxo+2F1JODbzZoNbUcxqD1z47f/1BcJUkztDUl73De/yVX
CNa+QJlMFDGIJw8Eq7bFOTwNl6rMqWNw2m/R7M/aBh1AtUJmZbZ/Ul1uBEEp3GI+19z8lakeMcr4
MJO+VZZWECVDj6kNvhCV67+l7Msl37c8OnPIuKqc4X0PsCEyJcMSCWkbbKw1Pptl7D9PuYFmZ3fy
gWtfv0MVPhjanLlb33kCbzyNWhmJGa8AXXlis9CDckBX+UgF3uIvflZHXoykqbCw5pKicEEYK38g
xkGhnN7qFnINM9J4QfqCZC5e6XVmCSsKSNH64cS4IegT9IMc3ZEZmAqQNBGHZUqGtsVioeejkrTC
0oiU13LdVNyjtygas2p/uhDJilBlqULcf7iQBOFn5TEOCB+Sg9qdxql5DMckCBpHhFQtcdmJ+fed
1uuj6dXqHIqvP8BjMDccAWklkbzirp5ZSv9aC6Tk3/9H5kOkIUhzWWObqMvif86nYsrioPWzoxIK
WlRilgKr87RdXXUFMVOfjCHviPmCrrwEl0B0m1KYxKH0vibTlunQlg60tLR+gm354/sb8J5oBYnW
78UpCmRcqfePT4rSJ5RWQr1tADnZdkE+ufMcT216HVJ8cZY5wVzQ//elsQCYNJHoslavxZJhf1Xc
4wUgiMfHz3k6qYPuhI+Ay8Xwcg9eoC27aSTsbh4qlwpfN8UWhr5qNdlcY/WZOlUn6FmkLJcFAEB7
Cw/O7ITNmm7u1+EAcGj5gapavoDqj492W6zvqHSF6DgTOoY7VQiyoVzPANZopBccai3ULOqC69AH
AXgnUNZvSo0oyjdXiNY6DMn6UMhwZoUwjbZJ4VoDGSIUyqgnSg5Ft5NxLyB59PuiktNBei3OU8jZ
pa3F1sBQOiI5f/Oa5ArNbGFvlOQry3dPMc6NDzf2/Rgi7jx2OA+kuk9BcKbskaFiwIEdFx+kqiPz
N6nC98lYcb/G13TfyQR/I4YwCf8v4N6BaK50hhNjGSHLCb0NR4VdXybQAT3jOr+sKWhX621VC7IY
0VwulOLeAZFpLnY0t70GTKo8/w+fZ3PI1kegE9KN0E413PfhimJKIiIC8IopTTRW0K98LBGoDKmq
Bp4/O9jyP97626CvI2u7oTiuNDggxj2ImV+Qx+/0EhXcG25PU+WQLXWahRJNL4Q0h0lertGrqcZx
fuczUPpnUhICxFBRbyABtJoVP80Syl/Rakbs0KUZ9PPsaedEEeWaDJvXRReJcccGvqBjS2s+7P4m
Nw0TAVR8+I6Juq8UaJBNASveqvqVhOjTSoeMbXwt44iVB+GYKyd7ByOlcyxDkmVJDfbwW0dsBBms
2IGUjvN8qehrp9yTiCoGDU//eM/MDxdWONC34SDMX7/+tQ6BM7Itp+wbzj1DXPHMVVZ3faTU7UT2
cxZHACX0cvNHzVPB408Pb0+0Gm59PvCxHtW4SM8wXmtlDJh8odydopBIyaGpxoQKUiPOhZ9NH+zg
At2OQ44PVuTC9jyrtzOr2/c8UlAuyt5ION1zU/DG18Xm8RAniaDEt/CmVbzQZ8Bs8pnH9TqQyUQA
PEl2fWgkAoiKrFsF2sGmpwdATcvrOE39RuDyqew+0zpt/lHLYG6vcWiZZvOJl3rCXYiWBp/B07BH
fpeD9GoraRN4BwlNzziPYIejT+uzzO3WFirpOMd3X+FHDMg8GflbvUdkCD6vkV0hsTY8AogQS1wx
26pTGdADiWSk+pi7OIBo5a9+KaJsIGvtnY8DmakMh0AD/BEnFU2Y+n8GbrFU52l/C5CmdRA9m8FN
3Lz+hFDgea+xsko6S2bu0uZAdCFvC9E+DiPsSAcGIppXttmCt7lKjLTz7rPgtu+jeRDcukLCvY4G
dBuzNPESsli8Z7OzbCZM7ej5J9r+87ikJie3L+tjFYwcNeooFMOxHLbaguFrl1gVFMvXOss5RiFq
mUs2JLxzRL2Y50ROmFiLjYdehq8vIJAMM6BgCzS0UW4qMBns90rnRME76wanbsZKk8v5Pt+C/I79
EhKE9thkvHxLwcjcv6bdV97d2sDJFVR9vRtsILAiXRiidblnzOuTXlYBLS+7xVrXdlH77cvwHFoF
iaV8y9j/5c7wEJ79LjkXkchfqa1LlAkGeegsbgige0B+PVVP6zAVv70H6NZKRPbhq4cPFOaolb/0
odBIvkWxi3lBYk9zGbrw9Qhz22zHQjmWyObMTLvHI2fXgfF/OHffyxxXfMTBH8kYoBQWK03DufU/
0kevC0mYDbmrdFh5zC6G6801p2hZ+iNTP1RIXEoq0Jxed3gD1lLLabElNMxAjrpLgZYiNngiFjZj
rBzaULj4i8hoTtGC9mG+ZUd9MwNZY12rnekXviAHdYcVaLJF7r4JOFO0n44O5Lii7A+KYMISBY3r
8y4lSdce67RodfERZaHhq5m9TrLSe46qfz32eKGsrS/TcW3XUKfkMQg3I2QVCx7pqgw82SLSVut4
+59mL+7jmohpw+CKNDDMt/CVKJP5m8Wh9Pm91Zij3KoMB31MmFsXEFhYvQ5nXwxNKOa1KkJ6Q0ia
PYKXIw0eAiUDc0w9Qa2tUc2XPrIKGKiY0Qcml+JEXaX5O0BY9lzA4FD7JXmuKI+Ij4fbyMYf81LW
bEoa4EmkP3OSm73KghZd9JLmLnu3osWBiVXdyDjunAtmDrrgrR1z19JXzfua2IqTl1p1baeclklW
ChXdTtLyS27nKay7dtZASNK84pKywK9q0Lc50KriEVpX3UDZDcCquFk957IhTH+KGMO2tcZke+75
Qm0Gw5xVNiRsJQRFhIh7wz+Cv6pTFcflkNIljzQiFxcf+5AgpckdBC0eYbyh/JLwx8OLegxzHj4c
6FxAE/KXCtdoE8MeriGUto9V9YSCbtd+33/WsZXgD5UZMw4Qnppt/zSo2sI2RDYgVrNfTopgXk0v
eU9MoIuFC34CcIQ1dQ/XPWt+sqetA979TbhXkAKaV2gFKAtoZp2AdNFsPXhfQxxyWFxmd3atys0f
JJpnxTgPDepcJoyNDRnOaERy3HNovvy1Kc2chwKP8y+A/XzUxntRnNd+stOqcBfVF1o3CEUPFq+P
zWyWsc4tZeN3WXsL9+tibwtxM6mpO/6q9Vmy+fV6hX/ZE1h4ped8lSaNProniPFxB3FO6gZcy2fp
lO+CCqSRHqCufSatktHMT4OkLxLkMJu2M2WpRlfc+whyQ2R0hT6dCbrI9zjGnmXjSZgKL9kTFfw9
xTJxL7b41KnRxzFolAIOrOpQuc77pooV7I5M1BSQvLTF8pOHhKwpMfNCXCce+L5LNZecE0uV1/UM
CDVjTp3bhu59HU0LgSt4OcLULrcpbK4gVpXBNbic9RIa1RVwk60aXOp/dUc1L5sUzF3szt8YCy+b
Ge+Ns+9cw8yLxS6c9tQo7KmOb5zkYKfG+iUaH7Dec51j3rWvgrRe0vyUYAk9ArQtTwybj0kOgmfh
cv/fUi4TGojBAS1BNpNg0fFeqsPbItDz0tI5cb1CbBtd7gyses9Hc/6PhlNrZ97Gcs2J/0U6RziT
xwnhUlHJF7TBrbE2jXScEOezsxa5Iw5m0TkisQudYnyiu5XzUksSrRRzsscRKSK+BnREgApx3WkN
fby0lSUUJsGOCUVNgdtV2pkNEn/lb9kSVD9ySiQJNsvsKUPURdIaJONueLkgOFiTT6lYVOzff9EZ
3IlZrsBHHhsblkvrImTbcpT7hpT+jXGvnPlVZONt/+e8Y01lPilYncl6olYz+rTj5xRi3Bke9zoF
CgPDI7DOL/nBFUgyqq+B8P/TBsYFxduHv/MWr5UHoFXWNcVYo4mcaxFPc7X6ztbz8Ea8KH8hQgcF
W5TnGxQSHnpDJs+ki6U2UuMiCbpBDakDxmFYa/JEI1ogaheomZxpI3t6CA+TJrOWQzW+9xZHc+Mv
bNwmwn7ZRs2kgRVhlvi2xp/+ZcSIE5xbUjRiNUfqpGwgKjCbYWk5EJ1rmsAzy7V11Mg0otFAwLfE
RbytEY4FNTLAFypilUl0n7zCg1fuFxFJ/FQ3XnPUA+2mehgL/rRdLBH4CGC7XVm2WK47xod06s+3
rtT3ltJMH9LLVaVWFRB4SWWu1rNjxNKU2tnrzfZI2jdk6pRGVhwgVYihZunrrhTKC4/kXvvRGBQs
kDU8Nyfwa7QIIp/CGUsi8ZG1O6aHyigQtGtXsBWndHGLYljH8Nm3+gQi94O4QEFHvLaWGTqZ31w9
4IamNzJdS7Bv+JZQJIp/1V3fiiNS7PRQ6Q+HDaWdUOKK4uhuESuYNd3EPWlL2pD0WIb0VtavPxj4
D8usdhBkBgnuHf8M/HXYSPjt+ip9oBlXYsJnVcBDR9te1nh05F6e4Mx0jWN0r/azz8OnWckXCcSP
WmDRsSTlu/oMHPNb38u/TmozL2+k2In9XJKSOo9B6Nz3paBS2P9jxnheBIdUAMzgzJDQCJpbSkfH
w4GLh3V/Epi4kF6CoSPBTbQF49A+jpz5fGpdn+hzplkoCeWaEhonGjQcRZvxFDVGTtGT6MtAU5GB
sW6Uml6GAOAn/YbY/+e6zEIDvgWgZuGkgxnzdBbiKD8NC/5yaH5Q2cPsqEDrimXKcnLEoWebpg14
k0t0/rAD/KrVzKfq8lQrJ+oPi6YGCsPDrZIjzVuwVFktg5OfmJrxR1K4QQADNVlyekt6DX1NIQOt
plGEQanfYJDcT8h5kaklzAl40UFoojuRGP4IBczhKceX3zhoNcKoDFbV9PUiDYlCDdQ7Rcc3BNT+
2stqqf+xHCTTMz3XOsmC1Rs/4sycfCgrq4ZmSlHZYQneI6tyJryAGy7ZjYclabaqpOomeWOpBGKj
TaT9OHQoVa7BkSEyh7Fw5b9jYTretMQpaIRWpURG+/QBT4WE5rLivCqYfWmPk433DHngBkN7iO5J
sLPlX1YhZOfwCL/lUAWkyRaTWup/KSFxAyHmYVtQGz/82JHKJrkUAZaQ7bXI+ONRf4+Lfj5Qd9QS
nuO90mZsPX+0aSs+fM1K4hNFPRLFmPzOJcRS2weF7iHjwiou53PJl9F8mEa9IC8ayaOgeMf4ckQc
c3HcvWoUcR4fw9zilJC41wnDnQnxe1gPHlbRIkreLMYARD5edOMmRqNLx8CoGllKPrXULf8P5oEQ
WLoras17kOYC9YL7n70G5zlLS8TepH/vPU/t6Pn6VDAI2U7Y7RQ2nv/X5MRDFpSuK0BW5Fwn+AV8
AHckvFPUsIbmSs61o0Jt1mfWMXohuX97j4nSdqi7umsBEC4OVH/tk6AKkx8e1qcXp+h7z5dNnprY
EomNhBLcKFdcoSSL4Xe5nynpEZhZ8kzrAyB+oq9mjogdakABMst/ufI0HPNmipHOK8kMFomNWlAd
1nGwm+gm13bCBKMGcgDgEiOXysV0sO6aue3TadK9IHL+opAvfB9AbgcHe96ZSDHOeolh+XWpGT9Z
LZnKQbESNImB0Q1RiPyt0xHJadeNzzqpwv46bqioGGuvDtNgeOZaTEgYoVvsEZykQgYW23fsw3EG
+8zSwz6PSIzTfoKsQjqy9qxtaZBB8t9+cxBVmqiQtSZeNE8PhYja5169IWrA4AM89hrWKkayiKYJ
SqxEDLuEr2GKvRx/Ww4it/ObDRX83cYagEY5/0gtL6gAb8RLVs+HwVZ3qcC2P/y6cHydfWZ3Vppx
FXOr4BSrZlujiud6P5iT5S4EHeVPz3BTHYrMUp6ZJCqFGdpHJEJciH9hSWIzfxSXbIWj5jM474ch
4H/2Bm2GWNath7CoWwePiM40mlJ4Vb6UeUrfaGpSQRo4hIUP8Y2rMHedbKWcRQ6ZbSYuHRi/Wh93
VH63/cNtyvOC0V2i2kq/a2hcSN/Bv3bQcGar7dkg82Hh19KW9syJSHfahtw/jOB7+islCGpBctsq
4KSX6epO0Nj3b3+xWgEGJIM/nawPDFl/VcCmN2T1yVPT0in3/TccCTMh0HPukxPCs4zJ26QoP/Ia
tAd1buOboA7isHmCYhGUb6tlcOlAZQ0OFEXeyGucWAN9WgfE8c4SU7+sSqKKwC/j/m/A81+lMuDN
7rWjLZ2f/sOVGxKoNMNP3ricQGd6oqAztfHw0oRDVKRKhQA2vuXrZJrmgD56RzpTcJ6gfkcEVjpR
JW/z/GqaZ27LXIY/H1Y+5s3PUXv2Tuthp6mD+OJ52rzYZHExOEgej2YRPNjMAa4xSJiHA3r64ca1
+Xccg1qN6RDQyHdjgaWQmGeX9ehp/4WiPoK9nqCL1AIKu6j1snBy888rXdD0az4zj4/uqWbKN0Yk
j1Xo69xCH2e/0mg64MtpBWQoI8i+cpDmTtCd6M5btiXzP8oe7iO2m9dtsMtZt4j2rTFcBGIbBeA3
gzW5+5GiMgmiy2yUeGqo9f4G2oxHxVWq3TeO5DqySO5DwmO8d8F53aoV47GJ1T0oN40PYKB2eaj+
dxpeTuQEqOPVvprfL/l0vOYz7zkPTOQrhPN5MOpZhUIL2QvZvfMZtKo11XTARwF8D+Abc3M53q4S
d84xB3NCZl7nPVG44QVFeGPh5fH0MG/4C7dEM6Jfjnhztfs2R6QgHLF+0+JJCTnjg0yCAVcMTi3+
Z4p6T5puhyDx2E4SksfsEt0X+FIUw0AsvatNFQIoHqEphy5QoUmgkyCZq0Ntfr3PVr1rxvhSDX0C
8eZLZ09OHYK4mYepy1671wOJf10XAUVby6nLYuOUt+gvq+8QHioVBUzzzA0CXDyWcJQ6SYAY4E4Y
CHl7N76KzAvf6UaHuvv9iK4bkqFQsxgZnjGmqrD4pX0wPCFCrOqVvb8e+u6Pe28rcj1ZiIV3bvpJ
Ex/lmgxnHhCzScjDaRSdVYCJ/gp/GdlouDQV/UlQSvz2Bmhtioc9aEZkTMEyZEAH8xcgVThIusPv
mY/rzTJIu5U3rMukcR5lHQaaxTRSuWiYxWJdsD95xH5XWXtEuRoOMRpmuu30EuiAxZs3jgGjcEjv
ccDPutL3BvnI1qrtX9QyDcX1NVXRekHBz3AndjpTeZHrKF+AIratAWu84H27ovF+EDOKGXTCwDnd
S1uMbmeQQxQELbdE/N3M2VfFP+lUP4gnMtFtNoiYGc3QKSY7IVgPwYk3lflzBuuvbJw0VVkpJoBx
HaIZCnkL8G4QakkOCv0hRNUPGfv2NcFJr6aNL/eaEaIv+NCTjv8QUqcP8Mq/i7IavuiAhI0+Udq8
fHhIWNMr209hU00eazRaEQ5dNYxK+UDu34BM1azPV0fTSpX9B9r+AJIu9EW7OJCoeKiMPUcNqsl+
6o4rLK0kGRxYXKjVFwad5NQEsBTirc5Ai7AhY5si8oiXCHypXL4LTzvMyhKXaV2qaR4HH7ZKHFdn
lPuBPxSWWkXd3ePyteT4fjyp5CDByZdVLaMFBZZ8gJYzjVzPn33lqUFUQThmyUF1YeBnTXQo/jwH
7dzVAqQnYoT1iOJJNL0SbDMhfRGvjwSusFzEmQlDxXg9yi0nwbTOcaCiJCY13LXUU8KyqTrEPw6p
i77H1GmoVRvmLUg3i5b0Kc7lFKsUrEWVin0b/rjxrXcC5vxPVLjwV/0zbMvDdLHFIV2P8mJMuAHq
7v+DDOJf9qJ8HWGN5hObS7rBjA1LGZfOhL04Y0jDOR5asvI9XqxkIWRIqYVsAgGzX/FdLyaS1Ysn
GsTaAekH1vG4D9RssZSYs9Bt0uxFnEHcbH9kM57O0fJzNboIuYeufh31GHhaM7CvQFRGYxBxhx5G
8eOgJWVceFknPs9oyHUFaWuCUSAwvZfJTtA3p72lvBwUxVu5CGcTqZZg8To+M9OSyGbo6N+JbcoH
1FjGypA1Udc/t5e8UM/gEj4Yc4dWfTzZeITiofPJ9T2cC4jkxmGr8JPZBh/NUqRcvIiSd0z7C3aV
HdJdiTpPPOo4SK3eurPhSBKd4+raBqeSzT8h6UWxEp1ra8Q9Ox7AV1RRVzPBaeCzqCXwCNHQPSt4
ccEWhME0zikpVdUL/bPcdoGLbRMsi95KoBYsRtcDL/5Kc69L/znWk1QtSCnlYMLTpCwhpJaJJfQE
6fIARM+j4kzvupzxD1kIy2RL+4+yxgwYB9Yj7scWDvoN9GZdKeylPHSYJ6Cp1tYJ9rCxDhEyibsF
7UKJz5m1FbsElW1d2ON8wDkK7SYlJZW0NlW+1KjWSAioTFXy+X1AfF5DfwBn0KzmOpWpSI3rJE8e
lWPGSuCGgWJ0CmQASG8rJ+gbREBFVVyOxzKuuYb4q3jojmvVPYeuAWlwWcUNNBAK/gL0FXFm6UYw
ZeCai/PZbYgeCAniC5/dB+lxrySSL7nvohR+Si8peRwHFlQI4JHi5NFWk7dAE4H07R1VwnIx88QX
7bEwZGxboyeJwZyZfOEH7G2UY3ML7jcLPS0tGo4ABGmRmCM21JFoeUj1jYb3fWF1BMoRCR7Hy92L
1PNN+2mGiDvmC21Gl9x9eqS0YbxhENjuWzB4FfzH5U9ciCxG8P38OjPD4AbDlZhDI72i3Q9Vh3J5
67Sa5pCb3KEdPLq4d97YuaRXhUI4JN4qj4b1rothfROJAbJC5HXMaety9z1HW6WnMuO0y/gesIPB
DFv7Fq4YOcujdNOUrgp6pdJwFq0phWV/1VZzndT83Htf8FAULX4dF3W1i0pBP+gKGx/mP0DkptrH
tKN0D0DNqdI2tkHJHfDSUdLw+TYBs0SW6vJBhUcSY994DGQUDfzeYiE+iYcRkdYyAZxL3s1DG8oW
dhjRwcmEZ0Bf3KGi5p12S2ym4kkvea9e3U6qYZ6vM+/CkZ6UWg5CrdTyoQKMLhKi7qEd3S4AifWU
kemy2Yz5yhaz8vomilGbeTrFI2XZpPnea1S3w4/JNvBh64QAP70BLkrohKn5ocbqNW4GCL3L1W0W
nsEAvitw+nxfqjcL+WCw9XdxiGNwKeX5B8hYo5IcnpBeNm+YfDRTa91DaZEFYegL1dVBHbzRrgae
eB7I0VvP1tRfnCjDt/VsIkTf4mfyJz6lfDJv02ixQaL4mAFwqPZRpxOcPcoCYQm0IF1vDzaiDnuu
90LB4Mfw+879z2U963FwMsXXmrPBlUoHis+xCbSXK0CEF6W7Pi2CM+bYO10d5uV1Jy7V1DZMfFHB
TSHhPBZ4z8/FuaXM9utA5TQqUKiVuL1iUY9gnKUwsjdUPw9R6284xakAKQrEcLebumNjGlMTBg7t
TGXfWjk6ipgVIZNS88t3u3xbBB0PNjd6HTEODVPzCDUdOriHDhMDAgQ8xNU3nGq64tNLVykhD4tF
WPhNaDQ0g5qxke5k2YZrlINrn5mwzQcsIx8aPzyZlOuz93D207eBlGRN4jo/OXCmfvdr9FhmC4Jt
39ACIzSg3QUWmo44QSczrt2tQD0pzGn8SEDYGFOperzUYXdFqfjPWY2HCsl7ZWnKGa/0IKTNX7e9
tT+YbtAQJvAGfjf8bJp5aJQx2AbRbDCW/ErwQlBpysIogZbg5Kr1fo57dwGbW3LfgOpctbdIVZn7
AtucjtNB4Q44aWBMj/KY+bXxoj4azfUrmMGxUZsyiNNNQqW7StCKfuEhoOfEYW0MbBEuGMrllVyp
6r0Tc3Z7O9HYUXv0agEMjQgpCsFrGrpueVebanUd0YuZ8OUteaErkMi+qeuUiaOX3SSFOMFlrD+T
BJyah3Tlq9C5JOObZoAbLrG+cQe6kF/jEVniKk7M985aCTHN6hMGpSdSjW2hctNtOIzD4vyixaAB
uP+lxYQNgx+iYShRhROB3CVF3IYoF9le/xwYrXnjNCrFFVfYRhbR8Yu3hH6XKdOK1FD/LOoYzBw9
iBnkgMDV4rlII609VMal87EY+1Uqp0MFVWYejqaZYwG2JHGO/6aavAJhNJi+gfFUw+j7cyLe87Om
8GCMLyFXM5RJ0Xi6sCIiuE877kaRUTxC5pUAZHhYDpc5rH4MtMaAffpGHI/KPnido6IjkxePBxh9
UNgLRdg53VsIXtLiNtlOQlpWm7xzBKQiczTiEbAozU74lSQysvUIA8j20tTTNNm4ibTCN8w63kN7
jiPMEC1EdCY7ktSK+6xzE1hbok/RmEcy/Sw6K5wlopY2Hhq0vHQqZNZHngHewyjJ09eaUzAotsdb
qHCh/0S6uw/Z3Vfpdeo5i5y5p6ThGcQs3hKxf7ma2XYLBn8IvEroiUsxxKVzXWZcrSkarQzpZFzc
WT5rV034uuFIYsSA4DI6EiDhqjVW+v29HfKo017IWMTitHfw7TD7F0NlZ+6mniBm1KNp0ox+FbUV
s0K0vmcEe0oqVdKY9w1PTbM5yf9d7941Pv7FJNVc8xowZlHtXt+oE2em+mBscphNRQgW0uGxB8H+
cnyLlsSmAsIXeeKqi3ghOFx6P+mM/qkAjTCWqHbt3cOdqxBnJMKxoqw0cOpZdQf58y/H/1WevVdV
Y+pOr1BoKtTXmBMOsEfDK8GBWlEgEkHpB7qPKCZvOPnFL+hK6pmw8d9TsMyw/lEMDa10Keql8XR6
vHrfxR+fXqFI7P31Oa4LZt8N8YEe7WvnLQ2ys/fj4+w42IESQ2nA4EeMWM0yC2JRk/nVRfGkbw8r
4XiE9K4hn2hDtyS4FsbcldliWFn1j2af5JiAexDxejcj7LiVviw34yabPXepEd4+C85VmUJOt0OS
B/529p8zkJ8pI94trwmembi/01BOUFTRkPuOH+OY3QZdsrY1wt+F01l4/narT1feW5+itqnKYcAx
MM4ODTH+IkBSTDow7HlNKASDladniIQSwUruR1bSegTQYE1S8b0xQc0gbFMF4hYgjOqVKPJG1u2/
rLMo5sjHpQ7pp+C9eW4g6R4xuvOvPNmyqSZcTGadENI59Bg9vL/6Y6U7d2KvANjAT+rFOdwnCMAO
QZQYJG/hlzbV5USylXK1bO2eTamlf7iJJ7PGKPw0qY1xHRfvAovt9bQlPwEZjB027CAdZZZPEJfW
pYtsUZQq44iGbLA3hAXyDYyswzUFNKqDOkjzmjcVl1q530xntO/elLNXonnVw3kOGqonJgIYMH3X
Hy/D1x2nP14ufsF7Q4S5Rj5T4XBLa5Ki0qqK6R+CszB7I6ROhvyJg9IDSwz5G81fRRP+uSP6EQTm
Abxx5JwUlNpuuQWKyJbiY+EVHMh/u12RwOpGi0ecS8jZalqo4RI+LaM3fcWWS4dpyux4C/pCkp0O
Y/JlPnLZT/FFxa5pwCvFkAKcizJSOpbEnXLnA/6v69T0eXRDacBIFpiXsc2OB5JdQMn9266fTwt9
ZJMWpvoX59DiP/rmX0Y5b+b2w+eZVR4NtSw7EO3GMHbQW/0W8TGcG5pcW7zMKch04HRjqPRrGa0C
DbquaMv3UHfFA9iSCMCs8cQruNMNG9cGB8wUKMhdKvvBPWhZehJ6CzjjGu2Bicvle+u7jiGR9gel
CfCPsF+S5PUyPCqNbdzowMDPgBZEhJG4ZujPyfMMDF6NIhaclssgiPh96bEh7mSXjVmYGKDQ5BZI
Vhl/JbSdEMXxxl02PUNmiSEDmRsIcUZzsT3e9XMoHRYDnqqmkiQbQAwV3zsrRr8lu3qmVM5iw/KE
YDXr6pHZ94WANJcMjNfg861wq3d2ed9sK6FrhM/bRA6sftWtDmoeolfJJAPb+BMCCsIxVg1VVl2x
dXNWZ4WCL7sh7E3nCLftAlMcuhszEPlUmlsw2fm+6Kj3GHlVLDFjBYrp4HmeyiiVVH7gWjOj3xsf
HVxGAIACICt88YcKcvYg3iDOZeymKzI/rqLuuQK52kvDepaRz2c/C+h7U5tRgpN/xFSZEleXdxIa
PA9b/DQQslJBhZXN7LHnSGdr50alaWbX5UEoM99KW3DptfKYxxrkmrX5TBy+7gmQ9wOFiCJ8awOa
KptzkVIaBRCfBtjpVeRNaifcVh4BpMSMYnwXkUnoAT6ZfPvw32H40/02Dku+KHqDqT+h8pyfmGY7
tlevumXwKDTJbNJxAsFdctlXx6+BPv2QIBTDUJU35ZDB8DG0IWOH0XKTf4YpMict/r2B4fOq+5xK
sfNNlx6RZUHXYvu54+Chco08em2XBlqaatp4NhtMdiILqUXUsasc1ecm4UfuaR0FgHGaFkqhGdMJ
t/t8m8ZYeVuZsS2sT09lryEDmfdQXcwdf4l6D/K18FyK7C2i5vFz8Dvd4UbfBv32reCLd7yNdNS1
AemsswyXXGGxKkx9edkP9Y6SetO5UdvT598YslNS0gb7vjC6Rjp7nOTC1PPjbVb/cKq8Va5fzevw
Uq/MQgeP1xqvGlqUSgcgAOW979pvbnlEilsIEv2FdIqegDfVlL2IIGVi0NfFVAtpsUbOFxtOOAYP
Pl+wjuEY5FkUxUx8HZySVb9aT5OT9ItlzVsoD9KvnqKXCb5/iGLerIQXJxgF0k2hI9B1ZMh585xB
5DwY1cXcvQHNuyV+t0e6FJ1yiRbOJ8WW1OQzFVkThZFu8HskPRzcXAh6hW1tx7dG6vKIlpzVxIR6
hUH6jNV2GJE8gcAPBW05SEKpIgjGrwLcKRphg5FDDnJVXhq4f+n4GifRhmn0M6/2APnlbwtVsBHB
nXW86McuJoXIOWi/nMicnaTgUC8Y2T8ahJWpJp1DU/0DfDpRon+7Pz4VJOD2ceX/nxJOmjiCq5ij
5/CMPINwjZNiWtAcUbP7977VNBnOEZauu50WA8w1ILZleHwxOyuArAg9CKKoBgFuvOAXVKvrqZ0U
6d1vWW2aZ3pQETQF61/ipO7PllJqo4ldfdn/e3rwzQpFu/ypnw5gAn9PqeTh92AOzAafnnw1PEUA
RJucFb4UD4BA5tKDinS0BdzBqOo9IV3KggT2v8HgpgUz8/E/JMmTm8Xkel2MIaVsfeM82bU3nwpP
g7Mcu66acGzB1hmPcaN8pkr7bfGk4VyX1ErEh5oJIv+WJgPqhFRkP4seNlrJUuyPVOeeSPvYFtNY
TbeEwtTobPz/cWAW19BW2fsrvDIDh7JhKJDiwJqgFD+N/jaufsvUmth9nNP3iHU4+7VZDCtjiQFK
bIKxuqgS7pc7ldbAVLEXCpYt+36Wumrd2MVc+3BwgXDO3U6M0MizZ8sQzZ4TlJ4OYvIE3eP7pq9u
poOxhMQBQqCELm5qAgyVo7dkGDALxNmRAwB/95cWfK55zO7EkpIFeCGjqMX/im6KbGatu0+zVUuW
02o7YQSGTVS8b14MNk6/aSnjT4M/+3noWTO0Ma9FBSMjln8hQZjhqJMYylZYwwqF/9W8hSNwhBiU
LmtcTcGUN0LGsqbMaTcx6EyZaD94WdUycJYSG9fkOHh8Ns85HcH+Uq4KF+tzp8UdsywEPab0oDVl
nKfV5F+/r9slrqtdueBhoqyjNvxCHBJaGGjP9OoxbGTF69q//5N6NmPi4GAGGS7scX25d6HGy4nG
u33kRVSXYGh9lj60YQwucsKa/xv93BO6YFWmN3Vb8f/xw6e+vxqZkX2PNCjAnjAnAyYuYKCFc8tc
JcYWu6s0HQu6nuzlqJH7lcGoU9wyGZjlEgwRce3AGAhktXkeF45a+ufHAVlCiFKnfcCHJivYxcQx
Mh/vTfbcFazFT/4kmVdIdLZ9MdeXT9L1YwpBqSmT7YiqpZM31CO/yrd3dPwnxt0ZG8ATA6g8Cdwd
0BOfIDRecrd2SAZu+rfUN0WdfTyprlFZqn4zDY/SZYPA5BYj57fpMslU0tr89qpFvi3mCFF/Pxm2
nk0f1Fte7dfXSdCqXSBgJ3Wt5PE3+XllunxPkM63z/JWLq3+01eE2VSbae/Ue23cJbHRY/CjvMoX
EAXsx2Z6Cok+38XELlbznzgGhd4Cv3ZYjVoNqG70m3jtdCrgd3wu2Zsq8Qoj1qwYRqevf7T0S9HM
tZsAjC/BqZuYho5WtrSbw4PI+3gS6RXaghDF05Ir+jEf+kxrUWjcjsQY6cP1gSEsVTJnxU8JdToe
o9TixF7tIpiRAYES+f2iyHz30EJOLoXvIy4Ct3ne7N9A6QeqPKsn04pTYRu1ojhiQcL25W39381J
/z7HeFG3UMw9SJyUsSQrq4z0wo6UH1tHYN0juZmlksHEqh0DtbgreeMbngcECadBQzwFVSxMqbnO
ei84sTFyBp7Yag4bUUdMEwHkpEb8ncrxw8ujfrj9hCkTtrPvD5K+B1FIBfggINxIZbcIL2AzrUq5
K5YjXK/4BQwTqDiaXjQyKHci/TGldr//OKIrCjt6XfYoJQMPD26++I/N9soNQqrdb9akdvEvEN9M
HV0N7o57MvHjE3gAi/TC9Igw8BBJ9eFEnncL6pvLt4066WXAgdd29VepyxGydp69KPN7VbwdbykX
TQ/MFejethUFzrthiGjQ/SsvwCrgowVEDkiWy/Er6SZrj9NYPwTtr9xC6eIzusbM5rd8Nvu/Ta+g
Tgxih62q5GrmPBtikvLvFZNzX/N5mmU8e1Wevq00C2VQpKo4VOHCetmuruqNnmAzoegPC9V4t+7A
h71k5TeL8VQpFYK8xHU0971CHhyWpXD63lMS2peNwASlOjdw65PAD6IqX6WaBUx6E/vr8mJntCA0
E62dcePsXd5dfVg3pWM/NdRiwPLntbrIjudwPEXEmF+JDzl8Q+LTx6TCNzQ+/aArwo4gJdVX2H+Q
GgkLx/nr246A0MEjO34mGZu5ni19tzL0U09WIgBSUzWoG+dXxHoyFpV4+6eGoTCn/HRFKSDfOc4J
5zC/Sb5UCT3fvRL5B0m+CuuE6mmpvCYZ2zK0Xf/BiFxNaGoGHooHn07CsF0NAJmmYJoKQ9RknX5c
Db5DJqXoY3rJqi1x2lHh2B9EVkznwpQ1vaUraJUg4v6xVIk9rBHn4Jg/D0pijx/C83OVqEx9vc+3
KfpQF7vFSQxsLz/UiZbKdkRsD0FuMXps9L6/AmEA/atmhIknl/XRRUVYJscpCpKhDxM8q110pDax
yF03H6JdqR3/hOKd4i/SNYOni5k2CxQbEhCYd+oC2PYdHCew3Fd8eAiD4ns8AqhRM3FCz3mha4cO
QR6sRyS/oC/vifLXFkQdF6n0wSVzR8A7GloqLvWn+b05K9fghFS9HBul5MxWse+JRihxgDV8cMAo
qMuOrRgitGdAxhxskTuxpUmdu71UewYk1uWVI/pAW8Hr9dl4utPC1M0gEm2BOUc43gOiv2Me3ZIr
rLqBih7LuQPg4d9QC315TkSHXl/06r1aAn9LajXk6J1NY9WANEyB01fkLUa661ojCjyFUJv9pQP8
lKFRdnOJREG0nyRgxX1kwoT8Ilu3k5t33v0MXPTDWdJc3h1mqA75VRcFR0cyXVdXQTl5KZe/Dlyp
5CwXJ8iI9Cwm77eqoRByQjwpFKuKxV6nZOk905gBNCI+RR+iKVFGgS0iuVI4k6zyPB8AHYR9AD5H
5xfNQpPqGsaBm08X3tbmh4EYXiuKOYG3n0EIiCht4E8nRCdfOqr8J9qlghTNiViUBCJ12MHbkb8m
wvZfjVVyMDWM+3DAuGKwCAZAUPFTtKSWCfMC0tWfqCOu8Hy0p6wv/Griu2h7QbktXV+pZt+ThQ+J
vn7+ZdMwG7OcndA27Km1Dsw1duYfMHDejMHMshbvGx39E0lOdkSsvGQByWOhOlbPoGOiPSEY3jEL
aeM0MgK17G8vT0nU3t0JktLbybyEvMYgqYzYNHy2jWul8K2IJ/c9R7jrQYT5EqumNSJ7rl4lFSop
lOubqND2fsv+NOYQQG18P6Pxzw5xBBfjizlwleWBx1XrFrT3eojXIjlxtedKDb7smdyt+COBNKtp
ixqrXAfH6MDu5zU0Zrd0XCLBuHSAQnigCKNDS2OYjUuKWBSB3GAM+1yInh8vuvK0AzzW0E/bPGC7
8xg1DS4w0SWPaEo5cEXJ03F8g+xPYCcIZmqL1Uidi9G0V53uw1q26KHpZexbG4EXZSWp1Q+4VAYP
Yj+5ytelZWOIAdDg97mzoqGVcGr1GQbLShlxq4rtZ5AznjK0EHa0FvSJ63erwIERcwhL9ivIjLm1
hl1ixI78r3CDxWAo42bEr8n3PgrdB2c89Kuy9tyjllqVUZ5/U+EKGNfXwDvdxMkxFJrPSMtLLTHv
MjZ5HnXUcloDljNHHDvkbxAoLOsmwrrKVUTl+DwbNsFaCRzjVETHIvVIbx6y2EHcCfxMwMpJeU1q
bvQ5sRYnkG+xpWo5PPUMKE+WtbotTRkh+qp2Tuxt6MboBuC7sPgaA8dO60XDgdBYTnv+yL8nufR9
hyVER4s6TUY25gUf2H3IAjq+daeoSbEtLKpBAgJEtNmHk5oDsvXePDZ+eARt9DntzDW/2dZMuTsB
Hn/DOTj82sGB2kPN/FsDrDm54aeknTOzbmDVXHiAGjZvGi+ZDF4ZnPwzncHVMAQYsVsJsMPO2zSa
O5CkO5E1dTuGKBx3IBl4TVb9RCGdnlAwWUhUGZDKnFWENXPZHVvJslOP/XY/JjQTrw7MDAt4DwVW
9NM/dkaJt3Hig0QFlDbIoblRYbXsdDceVD1JnI7L/018SLbLejMftCm+CXGlCzX9h07R0Y28rBkn
R1sURBMzz/jHR0cSjtUarlt3gfEVpqw9DMiuLEIpTvH1zeBQkcOr99PR/1umWj0aGs0ZMstEUlvN
nW13qaHO6s5C31AG2RzHuAPRXyIbWKtSdePZZErZq2ZWJafFGQ7E0xVQBO1ILAYuxNdNPadZ4hL5
EReUZ+EufN6yf5/pCBLbXBIaK44LrRzk93ajs5ozRHPt33nedQYSpduHTb2NOOW8mSWY7p8yCnDP
wUALi2kg2TIH+tDycAh9xH03+aYQm8Q0/kaJXv0bTwneXkjZb5G8KuXVDteIxFABcPBqLaXP38xh
1NXgICWPfj5MrqSr+2sFPkonbcpczfkDKgK0iLWFb0leVMFGd6CnigbF0eICSqw+IkqvvFMpZLD2
/Y1etg4bOoTWUFjKceyAvO5p0QSoiR3SeTGFxAhNLRj2yej7vlDSFG3uo6TmV31hULVO4mAsIgKt
gM4PKmZ3UfTI/rqIcV8ditinMycM9QTgh3chX3tWHwHKTI9cvFeSWgDh7ktMzIOB1V8LEifnkQ4P
6AsqRETqs3K3upsFVY23r1+Q6goxdtZmtsxSW7LVd+I6FVUsgVqlgK/DNy76tK/zFkYnPRe34iow
1bFqWIlsE0ERozOv9bFC795gi2g9vNqii3+I1QZR5M6hb+qBeJhrgdjJJWObusOzmCokNJxJafMg
SQZusZ/RW7P9e9vu0U9sbW7l3s5zSzkx7iZAAwoSTO7e9O23XYKX2fuA4TfErry6eyXHvV5v3IRl
rej/MjDSLJAL0fldqqps9uGy7vjOyFtJRjKpDsiBQuXhCam9mR40YSMPu2kWy35ED6kgaZYd4z0r
pcwB4H2JkVyaRhZkmXRZCMqBXDif7Sxu9RAJjzaZtFru46rPeoMF0LePLmeHGUNsB9L3wMOFR3NU
8VeibpalC6n5ECDGlyWfl/M2ELTuuzdcXqwklJBAbI+SDtEYcGHWlopaTn2WnxKYgyMjRpBzKA/6
8Hliph1Kohfvz0jtlsreQ2hqT/cyt+OEseU5djfB5lgRDuwMxoLNOhjpDzex+FSo31imXqXUFFnD
2oLgcpKDAhaHBBCfG2rkwIyR0TnU4nquruTQEhT0rONG4Wvp4qfIHyoxMqlp9eNDW1ywichXFolP
oOWlb1YVMoXG3cXOXJHugMiTfhbz21lqKHJyoTK19EPpbunq+A4fH899eyKMMSyVYF0tlkzuQeM/
y/56qM5K4qEdGhAUzC/Uz7BHUwRRVbCZ1cT6tDPK64PvkLJWHcrXUOqun7WyQUibV/gxsrhl14d/
Gl6SepWVv0OBH70GCrHZlH4Q7u4MXYwaLOL8pvwZrXHFYS+mnHfPjcC3KILQgeQ72qzNoG0u0fD3
mOuo7xFxU3lKTp98TvQRt00Nt+qVfbhfUtcEBvgZ1KJk2acwiMaduHSprZgwj7YZODd5IYKgQgU6
gsuSTlv2DtmaCFuypmfsHdCgxKx2Prz6wDNvfp8ReGOnIBdYym71lXjk/rN3mh9CaHA+rFx5eR3a
ZYR2SeZ+YoILUSzefQwxpJJKLuwX4hcvtfiN1QRFUxy29+uE/fsQk0vbxPiTxU/GKAJirGsajd0f
EX1CB134ZpUpgHy5jU3CHt29X4ttJ75mDRRMhYU9a4U6ZXvtNuhL5JY8rtzH++QIWrTFl5rGC9uX
qz6RU5bU9SD3cCPCr0E2QR312V2ndnkyzyEgdA40lphVVjOTzfwxs+wHhHuHdL7X9hzVxLI/TGGk
Ylds8oxHO+yVPKeTYwJRlDAzoMXw2isoUpgShMFhb26tfWrP3M1pMjCFYBwKk3fUdoOOkYA/fvHz
zn20C5lg3Io1tGP4PVAu4h9C784FwXcW9ZGMUt3ZnY7N3syyAh/9zWwNGZBNpv4qT+bBLHSe85yL
v2I31gaSz7Ecdo3wv0krmlrjT5E2XAXwJn2zHvCxb3j/5VrKUJI1YxOmr8/S9EqoqXOJSucvTG+Z
CtmSNWLh6p+8vxNU9MTYP54zehVzrUILqk3BF6QukBnwEPeuwvm/X8wQQqZDev7G1ri5yMXaI/Qz
z0n+5/qlKM9wt/sThPi/EIzjC8ghFMKWZY0NDH6zJcC6e+hthT783A4fLQ49okZv07Nv/kDZWSuN
UNs0NgkWIPhRYaAcyr7pjF993swSdFHtqO6rV2OVs/uCGafZ8RIuCEL8QGT8fWvYPiddcfGzw1QV
8pkJZrQxZW6QOOvBEpdCETNARf8hitZozk1Ma0K4Lqhv7qzAMU/FGWnQeT3pS2EnD3POjN1Lg2dz
8v85E2Xrw2uPW4c6oqYEkJISYGMgRj3g1AgTsINTSDHr3FV5th2eO2gW5KQebv/vw+CZDbsKwpbv
AvAeXY05NROqDDbAgV7iiM6SoSLgiGy+zd8aoq+Qw0n4bnGGocZbZaz3E3kdOYHSnbmCrvBoCh1H
SLEl4W9y/9VMfGP7HxunFAXrcb3q7MS/bHEDfp4V44Bbto6DfDgvXQlnv4Ywr2KDeMFvzIl3V6AU
zFJdDSZBLkGXYmGFqp81CmHu6cQ++6fJXmS8BZ/2J2/AK/X34o6fSgRTpDqyBWi+v43hGu9MjVsh
/KFu7zYssgOqMsqLUDDDThVKYUL81k90Y1EexROFfzZB5xXpPUmIttyjurS/nYyaVKR2PXy7k2om
shFGXCRThmnq4kthu1bLLQ1O5Cf++nDWV0ZhNyzHL1qEFlkdlr+8l0tl9C3uaGPJjiWXrgjk0ERZ
Md3T/N24WGppup4GhbLwW74jQp0FNbCdsVXIekxMDXZg5BnhDF+k0CJwFD9QevOyX4kHZOrFK8TF
Bbl/hkEqNApVai2OmfmXEO9YTUofdxkuNdF8xFpdJ/6QX+uxoG1ypiT0/NKJVg8HBGH3dH3vBLeg
UREijyyrGRIu+knr1bYWrqAjbupT/o59gZy+1e43/u+9wQO9FjK4gegs0BG/HJOfDE9n8QT4+I/+
Urkkpvhkh9htazB13bEUJ5JX4LqoSh3XkhxFQ/wEJmEyTDbNbi9hE0rJTgigrNeSoHrrQI1LJxyP
4heixq8Ukjyu0zuxv5a9YNoKu2J9UZ0AdqMopLUugDp7KcL67D056DvWF0Blplr/PnP8S8siWQlg
LKx+uxbl6poJvIXhGjWHtO2+zzcTHrSlnFFrxYnaT7phNuN5XP4n/Be1I5jhr2Ix5RmG1Ihxg1nN
p9PdbqEYF4aOrJF6zolSWOsr64MJg1PNOx8OndfnggjIFnBobN4DJPRsYUvIdKk/e+gaO4faGGBS
LGShtBBRLdWcwySs5EHhZZloIT5tG/vIxjjvTg9ybXxaYF3IBmcthptCxEJAbLSnUTDSvCbSeH5j
85icR2pp7rbj81DRiQwiyI1haImzJnGFcUMUb06G1D0++eUkwD5eqEtxsfQCwiQdUFr+iLZeejgO
6N+As36I3enYBJyzvy0BuY8xv4Ism8GiF9jFZJMXqVdAXgDQp5ZEd0fwSSLMSXVre7+d9E+VcA1V
BnvGyhGY7+adsxkAHIQmMMc1Np5q+ZXIhipwPTDoe3vOMB9yglHs+3byLN8zcIcqRY9hyMcwgJI2
uWAyvbbj981px2tJNUJ0ikSYKeFCkZKyyvwfJKb0h6cyN94KUMzGwJefUF98PTUE1Ua6lGPwsxKt
Yl48GvxZ3lET+SeMeqN1mJVR+XVP761EwADYgPl2vj0K6kCWb/0wH7VIJsKgtO8GpRNl/f5Ihn4I
EhXt8T4RIpT28j8VruWQGU1a2AHjxpUQjxY83TrJMX2qFk1tS6Fq6qDqDxCdAPCgrOXO/A1AYGUx
ZJCxkjIUwT8qhC5j09hjpTffDLkUEqoraPYKGcy2h9hzZQO817zaTmjpLra3XkFeBnVpXFEFjW3R
5aGdUBOEDmxg/IkKVYTGeta5Hj/qdT9bi590IXTm7G7e6VdImmJlbuQUE/fb56zYdIwlFecIuYa/
Mr6lUrTFCOZfgVbT9yuawGayu0Yb6gObJF9YUNg/eN+7RwqrWOUZf4AdCUiVFJxEV3tQRFAepmrm
UTjFrJMiQ01U+wnzgCZtbqLqLGZoG2Mq7ClKvWhoJ9aAcj17HpM54rrXNQ3k5fua+/BsnZe7vy3A
htro9xCjmJXCXqLWwTxIYeD1nmD5iG/m7Uk+1IkZ31UPiGz+H1cYu6TwaoJs/+uIylt6OXph55mc
gFpkZ9MYUsQzyBTj6DOXoA9Sb6iYxTKVwRVb/Yw672OHfeSkFAgz/FOxHkkWqeqkbPe4A6f5WP5l
UAO0iRvSxLZTC+v9UTVeKsQYzEQpp8a4AtNP7PExogcXsB7tAvvjk3Mzh7yL2KjxzHpzHrJvUKuq
O0dI+Es/tbphAMTlXcUvLrH/5jWO/UNFybcOrtDpDE6voyADTYLJhmHVNsgXyOC44FEBru6d7Tf3
Hel4LveQWwQeDWdDSgJ95wakGPtoIM6OgHjtflXdosFfWzlr6uJ0bw3UhThv9eNIbwA5WrYWdHca
WCgTIn+Hh5klU+LLmCjq2WBpFDUDSLz4TKez1QxWLQbXYUtp8evAsGaMvoALK8HGjplGX3CeLGdR
LnuIe+wpYaQ2EMWmeEBg28Igd/UjxDofA9BFSvUdbiSOhus8NHuiZ4Bladh7hbh+OOVTwr/VoPGX
3GDhnTnRhdn2TSHoSOAbbkwjZP9uLeP23beTPw+jREh+fmpmmVjQ484bQ2ve/pl3ADWRupxLbloc
jKHDL4fMIygAIeAHeF4hM0DexSByYHLOipo/CWFG5umd1igZOF5whxYX9y037/4KzIZrxUDJtEcI
3846GoSJin3lb4wbJwS48X2wAOu0OvBeOXEb+hXXm4BnwwbhZVZ4SsFLBsOZBzpuxGYnUngO5RJU
A/noze8YPY84zv1yMkJk/4kh9ns05RLDAsJpekgP0wLJ1L2bL2kW8vp3Hhnqkx7jz+AUfcUsrBeZ
y44I88oSXS1cKAnLLK6JPQH9fsxAStcU2mZGI7ZCSKU4x8K7i30f2un/ZawAojWc3ZRRHC2/3qXy
48O64hWA7ks3PbhjeXAh9y+iFSjqoAGNidGnlKe8JkWVDdt/3G0D84lBvbh4MeDtwlK8ckLRsbrh
bofUkQL7iCOFhW7H/Hsp93MFvr55tJa/qoF1iXnNxEIODW5J3uq9qMn+HDp2i85wECxiGqExgnEM
EZB6rhQzFAqTGne4pD8f7hkf+ywWNk3yZ74S+o4GhbYKUPySoqW+gJ7iArgfs8aVt/LZgyXD7fd/
nsqaNU95CaETG8L7Y8kjVxtg9d5EInQtrr6Vh/gmHp5vC5lvY/umBl0q3LvPcXEqKzwouZst4UVh
6NFkmG2CfYH5+fFKZN4iwYgdlJFC1JVolqQcKAMqYHB6GMe/1pFVfCJIYTbUo20mOeeAyxvXyLAM
2D+icMys+OahbXxcWi2J7UbbYcoGFdgZLhLOyMqxwdmWuHyZJAjZsECfVP1QPG/JWKyBQF0+YZ49
n0TkVajb8e7Q2AgakzryBNHB0LGp8gPMMGxyOYhx3GOgwDZ4tUkkjxCDbUN+GZ/ccNzofzykoSyT
ufO9QMCWbZ1Zd6mFKFjyQUHdFtWU3WjJSv/Q7VEbY43vNo1RGoVplWhyaIiiVblNZUgps/vCdBJv
5x5dgrOk3u/7uz2YMb4fnoE4PJ4KahSrfF02xyXG1EmynChmMIRr0xYREBX1I91k0Fb4PYb9IYm1
j5ZjMnpQYP2kBueQ/SneABi9X3Kf+D693Q0tPSoq83VEVIjDFjOWNQ9rCD6KYxXYqKauNx2S6Eao
MPxd3t635x8MJTu5/x1iVwU1J4RASJTcrZR6cJage8H7wEr8JnuE67d+Stn93whSLG0LjkO4fn6+
EARnIFdr+9pYxooIAnNxN8FiZGTyQYYNyGVPe1VLMSpq29ae4+DMap/rXSdbu8VKJ1qSmjRs4CAh
iW3aXFqtzCW9S5x4YCk6mk+eJ6nr6KXcJ7j5Aken1bCtx4C+Bhf+DgEvd4U3mX1KQeGf5NJ6Rf1X
+D/LFHnifg6j3MUpWEKSfQZ6yhQVb5WUijCxsB/tpKP/aV4BSVzgG6KCpmHx+VoSnrWo4649LaFp
8iHRA7jqTa+oZ7sj7p+2gi8C4CqO/YoiaqK7XUovirlJzQPumoc5Cihq2OR3Uy9t4QK4OfJt6enQ
UQSSghSk/Xci5+05GvOq1Czjc+P8KFNvN2dXNrGltmoAKAabSEVziouH2CewRnKBcleGBSJnwK83
AYo3ulUULN44ml+xTM9+kdG/ZHU11gwfA3ZyLulL3Rr4SQK1DDU1IIb7L0EALubUnpgq3iHWa+5J
PdQ+SJYrk18OyQSf8x2nlmC9pZ5vrtpDyx8/036AzsNxinVnukFpfpvnfUQnz2XcHW82ltN2SRJ0
GhHfmq8nq0l02j7MRdqC+VtgOXMN6KBZsSq4ayNYCdFCK8Gs3cahSKMkyQYdI2J7n0FczNqLFGK1
eBg4qzQ7n4Rx3sotRTyVzHXLdDXB+XCwKyTg19vPini5Bcqqd7mIpr2yAV2G2NDEFiA6ikRUWbWY
7wtCdzJrtCNXw9Ut/W2TRMo2bIooNSTM4M44PNR4AQP4CcnzeH4+WFr7sKf9u5UZZyAM0JXylLFv
wGmZle2xAskzSaLTDWN76/3TGj0uNeALrTXnYN6dthXjypovxbl0JnWGnJxuvf2KzXyKEJbuizKn
WIxWPyLwJ6hLCCXSSZmwmhTZXjfY1kHWKdUNyM6oF6F+b3iw2MbEWoFproGQo9QokST2i/MY5k3W
CPMPtr8j9OhWD1u9Bx93YcAMMj6NxxZVRMNjrPSxObd7frW7Qi1PaLmW8pAoFoqr9ry9y4E3AlkA
wH1KghPlpdI/mmsUkLvGC3mVZdMnHua+3s5OW2oitxhb8lk5BQ8SR7gwgE2T81kq2l917+hOuHIw
XEwba4PoP7jXDJqmSHq8AJn8AoLkqKyOS8fBjIF7Wmbu6zRPSLeViURNvDMAgVo8JvorPpMskacd
wPVf+pQJcoLn2R/dsEWAu5t/I5mqrjSkg/KBuyHkGgggPOfHBLy6Mab1+I3Qd3oreSDlYxWqfYm+
ii6OsEJT+0pDO/GdNPWFFIjjK/s1VhFhdb9olfJfyMmehy+lDuCrAk3S6KzlQX+oI9pTccE9Y3vk
t8CXa78szcZtRn7ACmhHLFPRJ4tK7LNC+Xa/MxgCSDovwETEMPNbUv+CfJiWDtMZg0OtZVltcEL7
dAyo8ZwLF7WoYoGKWQw078d4jss0z3xBlbvgGbQOW5XTLARlm7HonsezCaXUbnDuxe6suPPNeBqz
+Xh4vVZNClm7w+W1vc70yRsSXVmfQZigyAcuChBS6dOlC6ELwPkiz/OwaBrO/R2AQ1bpkGRShqc5
4r+naIgco4dRwMLfyok2iR4/+pglDQCcrVktjKm5zV9422e7mTWLjI6G9pODVgszh8KfplciZ0kB
vXJutizM3RUhiONYdaLq6JQUEefZ0bNI215BI/ghkU+5rSMfATjIm0hcmJapYvbzN0/3nlU50Lb7
3sp/y4v6pD14ItWLKX+Od42b2V14UdR24gIMP24eQkMCQs971IWf7jXyyvxg1QWitQKc69wZs9TL
f+BBwpyLCTtulpvQrybY6/ccEF0RUn/rZqcOW24eNsiOo/Dm2XBhG6MJX02R7WrsaIk1vHl/4lhB
/OffZVQvMTC88elOhgNFzdoPdXlHhVl2UHOBdUx8oKSkIa8p2t+k54UdhPrTarbuVty6FV09Amra
Aa76LNhU/gEDCR65cZ7CCSZpkzk1eMQgXZytyygrWZ/CHfDP63jUdHo0GZFYayyj8MKQkLRw9Mit
7p+udfPdBBM7yYGCMg2fCe96ZPqpo9dv8u5Iz5hvDdLr8CuX/bBWsTLvw7+9oBda3s/UnV+WZ/Zc
Y4FMyPxlLS5P49ucBy++dAOpE/UfMGA1zBBXMZsp8IL2Tf9TsU9wbxHSUhO+UV79E56iNNEoXv4f
dmjriv/g8fq8k/g+jpYnDFvc0r39X0J2BkbePeMkJzmNheFy5pgAASgGLAthspC6vXXAvFH3YD5U
sHwDEK3SqT1EdWvjs/xGuRdQ+1TcaVr6Qn+G6sSCyF30xo5aXgmPvf3oB10KJJj4nIXNqXQ0fJmm
dSvH6olL9G+f0Gxzcpfg9TB5rpOZ69OUbF61hB6WIKGrmqaGUvZgbh87ziGdNT10IGlWDhfyjVuv
6QEIWztgh72LpYVYEtC0KTFBmYHfFuui8Wu0iZs6Z7c1C5yLAYA0/UJwkuF/gp1M2NtJnSCzqxpc
v+UcmID+67QpZNFZUpy4JXLlaSS9y0AmffSYEWm6ikjiYiMKvQZzUJJ/YRpQjE8aT0/VpKlzyK2V
Hx7Xcvcu0uW3sr4qrjSvNf0nCtmmy9Q2YqtwKjqX9gx4LfxXnmm48GZNqbC0zFRfoz0fCgq4RqX6
S/93kuqHcody9ffm9FMYlcPvwDFOLYL/79USn5Ee0/PnfVgTOGiM9cqjPNKzpMrsCgcjbIESgra5
+pT88fnlsFedx7FJpw18F0fKL0oqSTL+cfvYQMJ+YS0g0ASka3EvTfm3Hx3+RWDHQdueRmK4nRL9
l3AuBC55ZB+6clOabSXTMJXTCktgFBYDNJtjbYhjDap2HwCLeOqT4jjj2I1jcrcio1qy+2lt9GRV
k4/iIbXa6wFo5xpzpp4EcCpGXzikKDlYOuHP6iwdwbsYpd7Z37TCoFvZ/xfSR2VPnyLTSsK/9fWz
6GhQn2F7T4oKcXWWm+ELnU//DVP3WvpfHaAHSxMzW8gl/RqtU8FTgu0c2k8GcwwV1dhn66SV4we7
YMk5+K46lNnUvUfa6HclX3gFWx7eZ6KXcpl/3sib7EFbSFJz6DKG1A5+pHRQ/KY9u0dlifYghK4y
Ap7oX48hQtw2mZwxejdj0vi+XCcagFYotHXXYlfyl06W9e6bdrcOoRUsug3t0b06Wy15CHGDrImF
3tqdmG9rxKi7LGNoGiSd+IKf58v8brjKg5RDN9yEgh4sgf/dIb4u1Sr3L1UcO7p96KivtQoQpHBF
i78IxQxgMkQ+nMsIB8TyHT8uZ0K+xECzqqZph6EGHVuL6zFQ6bzVdgeNRvRO0M0BDlfZdfZbtAbU
npDLNYvcNLiFzRdjnhXnWVV3byAxG2TyZHeBpY6g9rl00dK64Y/iEBZsj3iJqkX8+33nuyQPeCGl
+LErYanIbf9mNe4ubbXrgKNS8bU/Tdc8oKc9XwHQrj5cyyxiEl9J64OiGsG095O01lesgaedJWQ1
7FCkMV+nd93/eXoKaUgL6qoBPnpTlJkt1EzetlCCjQaFP1IHUe3bzeABhAOV0eWz4H5gGJa23bHs
NM5LU15kRpfj3NWUGmpl2Jn1/WqAPeu03zEibd2d/qjUgzympoMDdxtoyyj+6qnUU/v/zwWaE1W3
hxje7Fftqm31U8ZOpdUyMXF1fgae0zZiGHv4m/V0plIfne7RBPlMcUJsX5/Zmuf3FqDlXz15h4NO
Fs+jKLXMO4Owx9pDgYr1qy8MnqNPK9M1LaV1DwRQ6fKr3s40GpzYR1PvD6krBfzJnP8FwJngup8g
4QgiiZ4PGPbNkPAbKCWVAQccP/fpoPyJKfBaVGTUPAktTO38t7syb3LhO/dgR120ipuhSP1KRul7
7ADtuyvwLuYamnq5NXTNbSdhx3szaXeTJRPF3vQawPkHe8LUve5dPVFHZj/kgJy9Fl48+USP8DC8
YTuo4+nkb6Rh1vMUvdsffPiHMS+kINuA5xjg+fU2NFVfoO4RFOp5eCoWlP13O9c5lWxo5SwAka+H
IjS++P+Dsz5UOCAf5dnFGjXyE43I+KaYJ/pl5ey9wGRVPXDd3pAsSZsS1SxtvpE7Fm5pG9dADKEP
GJgtpNNPcSr3msXX/mNDV/p0sPwTou6cwxrqF1vlvAx/fvFyEM2CAOYVLIL+qw4TM9S9+1QRU/HJ
9CHw+ow5r28tH8jB/oUcOBtBfTqlhXp7CJqzE7dkfHV/fYrVRv/+ZNSIq2oSLsNFD2dC+tyTv11P
+fUSqQkWLsyHKGER7mILuLPYPV6tPESu7EDhxNhEtpkGmbu5HNntdKZB5v9YJeJ6FRHle6+HSfr9
FVSWwLA6auLmPtOCBz3i1wtPzLwasQx7V7AN5wXLVSHm/MQ5p99hn0xdNt8pu+51HhQcvGWQFzUx
lj/h91grMqZbGm1gHWffnO7VDvjtW9zuM5RsvsPrm/y9EUggb9H7TIGiDIPUlhdmAMvX6shSwb/v
ejZb4Z7PC07PpVj5dwsuTJ+svDQxfpU4zduBIWqb855tFUZYmYJvLsbtmocpOViENi2gjZ0jjaLu
r4lcVE90GO0b51QnfMyzfBK6bb/YbxgNcUA3RUSP3VJq8R0DAkbEDbIWD6iDbWxP1NVS4xsWSnhC
YAZYIYQ0efoyBJH56wZ/lqlHofGjVQ+JcHB+VIeWSE/m3Z6eST3z7cm+0eJN/2WpVchBgsSqLW6T
FlffU6XcH5KoRSl+CNhSFl4uww8yTtEItk4Lf8mSZJQGjZwbccp+uKs4lZg02H7/xbC4Q8yYHVT7
ZUttSdUr7Zn7wQg4pw2Qs6c4qBVWIMJL+iRiwmfGGAmQI5PtHyQBxaPIdjLaAtwvnezj1KtxekuB
pVMn8t23N/3nropwLW7rSSqemoIe0kmdG5QP0I85HWdTHo0ZpeNP+7q3FFNcAYEq68/W2onH9NHV
z0Z2kq0n1d/6DonbVp9MSVDpFiQdedp8IYMC+IO8HiP3essMaTX5JBR77QwLbZxRf/4AkEh5XnO0
G5gRPI9+dXV12SNVUzH7VN4RZDa2eIlLl5E5dBG0MRm6cUiq0uYymozuSNCbtPQjA//5zGqubB0t
jy8NliqDPZtLsOWiIDiUChkz+XIToaW+rWPD5lSxREuWCgeDKOeL3EVrVMLC1b7HGRk51A7jLXh/
03zkKPRN8o5h1NlB5VMUqemzSvchzn9B7W6yFaD4iQZsWLfUNFybOqWAOCGPZnH5P5Abm/LNPslD
SJb9KcyXf8bVoDQ5fvxixr5R7orYCaqhkwMqrYyrN7MUWGSjMxnpKKKXAsnu8R8rcoDtrKeUs3MH
HL3qlbeGLJPPxO6BmVzIVIdFcVn6jzYKujjJyE9CBT87/Fb4AuEjF/Rng3q5zOEZJ7y0EloZmpvI
JLSrSjtAQXBNpmxfcm77xG3HLQmwasey4hVba5ViiOsmdPUXbLufxBrfYDH81comNzY72xY87A3v
MricSeq9Z1dWdDdImpifuMJJO3FpoIv2LejL2smNBlcvNILceXXAXi4qQLMZJ72X4aQhyb7GD8/A
xKfJws9Et1H/TUOnwWhy8tvOHQqG5Q5+8Be2VvJr7BuBhR2eiPs6NI2OWDXVxp/lQbhWvRPW3k2P
0tW3OtsXzRkj+7oCaUPCkU7HjbEreCEdTPysJYaNGdwZCeNNCDI+p/Gu7aUtofi2HzKykzkGzhmJ
gyMDtJmC72WwaQFahSn9/IMEnq5EOfCV/+4UpBMhth3xf1G5l7XXCTVlyigPWyIiwhtmxQvpdHC4
esZ5OwQ7J13CgCBTlfHV78JXLSpbBAkSCpNcFZPnLrm9Z15jYQBxRkm4/HH5YVTk9qcij2RvFefn
FlRsLyTJkPl/SYqRmas0gS8XHZgv6iYMf4HGFvweArYvcTFaF6iQbhwWO4AILtyBkUYfz+mXSyYJ
aO+7ZKOpFKMuP//4tgZCa8WkfIGbv4wJGyTimGiG7qpUln/b7tt/uC4Zz4WS2prWWbbH3roVmAHG
hQ50oHTBVd3O9ekVBk02fmDcJ9bDCgDFOdQ4jEoCIsuzgsWXahZ0nucNx6iKEsG0cDOy8fJHwXke
gB/UP4xkCi3zp4KlUdQjf3KSOgZk4KiVU3Hpc/P2nEmG4LpBR/bIp7UP1OLdIXbDySbv0msaKuba
VbPfmBcIjfm1FShoriO5ASZojQvMAVNq2mrnwEEIkBjhvj3VfzFAV8sbFEXlKfMWjy66SGBBRZqA
KJbh/AheFKrOQh1r2h62h5Oi0jUNUau84+TUb35Wb2WjNFiCzpJk8eG8coPpWaj6iMwkjMaRhEBF
u+xQX3GCx+dmpNaou9I6jm/vUVQiTnxgTiDuBz0hnhNhRaUNUhscMxr9tGdJFeI9u0MSfMGiGQOX
/NC8LAVovCWcepbEso0/h2efUrpFXnWdRw1N/Fei7XilPp09WMGq1tGvV8XoyUEIE6BTZaA/c8iC
m7++wBUqzPszC/EbrOozxVSruWELLj03cVPUZOizH7/Iqm5MtBzNRGFuvKRowLHfnYUQlqPbEojn
I+nLOUFzzuZxyWRgvqUZyJ/ii8cZZVcejOfiFoyV2OpYOE3wWT9G0Ku8DuG03YAsYfIsn8CSvhHV
HWlPC52czGt7/aNPled7HA6O0DiwcciOHeb2TVuO3Hol+uGxaIQ5vGHqM/c2V/IEyut4/idxPd5n
Aw9t1ZTQaGLeLsxr43VIPylc9p/urh5OTBdaCnKEtIKmedPXn19a2W5lCjeSN7p+iVIGEcctYZ1s
0hoiIyRjSH/du7CGU+6y3R1AXUwTIdkAxAk+ZEmkN2pWLUnsrGtiuKaS1lAJvE0rxSAO+nZe897R
g5lW6uVv6pylYbnUxFoxj30LT82t6sYSLhF8yrYx1ytq1TU/18JP5Rrb0QE75ymro3uLLVmE8rCi
NpwaTMTROoYePIP9oX5m0bgVF9ORYSU8XKeljJ4TRUYO9oypWo9ixnbbZDP6q7qHMFqCcfK8K1cM
auCBFfaPz7zlrCGCBgWigDbCIgkcx5A+UtcJJfxpL0B9HpTwzo0TjuXgpe3jBtb8dXt3v6FKT8VH
HZwYzS+yhfb1Yl8+Q1p9oNff8tcoyAHlFXc9FeOwIsd9Y+B1kSrs85kSLNOhohnyGdJUwwoRk7EC
vRK3yNemOP+5UufWdcXH9G8jhVkAzP8mXNLJmPPrZsD5B2o12IyLQq1tddDmml+T5jK3ddoBw5Jc
/9t4SdnKbCz9rU2pCCZMgu1OWH9J3q/NH8GsTjqMaWPJpDUn7xKLTQTzDY9pDxPw/sDiwU+efzGp
1jDvY83ja+KQdKmJBg11+diF8X7wx86DpJXdZSEySb3wRMTAlY1zFZ8JfSjdwyWvoTeWAOyTb4Pa
JrBLb81/Ke75GJidys+OAB18LuWEDHQ4bVMjNTZUOTCZltojvVx5zKMJ+flII8O1wCabpYZO3GHa
/JMJSc9s1NNOwH9Tu4ndpIt8Uu8SLdpOyJoFNFmH7sP58s1dgM67FHbaSgcDheMG20ktyNf97i31
8iH33H6fN2FH8ubYYtuRvC+CvsiduOCxP81fVt9iw4Va/nZDlU8bnU88GIQawofkZqrF1RJrTsGH
/f38Z5xuKr4XBUF7+MBzJEr5rfj8niwN7B7+IrkI0Vv0Ed7Schnm+WVt8qr30XZ5F61SdCSKVAS9
tetlJY/fIDeChZDMRUT3Kcu51sOKfLzw4p1hT8F9SA9qC4Po1VyI3HSvwlY9EP3QLAOw1cVVxqNd
bTfz7VzclG6g9Ev8G/uST4Ia73PMohNugDz1KOGBy6Ydbsn/YT1eHRuunMn3cJVSz4vOEce0kNiB
K9H1UhRhET235WQwF/zvw1lVj8hz81jaXkzZhqY0mHZKItkwOFD0iwHAZGCTuYhZQrIOtNWsZsLs
pe+f8IWK5hbveekpLS47F5DoNIO8TD2JS8bvW8BYoSwcGi1oVvJvQv51EoCW89AQYZg7q6pZSSC7
p9FWvMAiy3CfgdXZc4uXRDxyYObOwo2r+85dg1orUlkNx8nJImD0z3KrlaC9T78SKBBk9BU27EeV
/kbVtez3u7qb1aknUq6ZNtcdmoxbawZ9inXyGbzDw53/ckq8zs4eOXbW0bOluB1XYa7smzmJBGM6
vb6wyLH5ADbuVxTlWC9iYDkSmTxySBJEwRiwQko888sH3chMd4PSFrtKD0WEIkoVVHtgbh1C0TIT
fQWhNRNtUgXcaLdyFkB2SeMzswejtPVER9KJlWOZ+Maqri5jZ6SeW+bgJJa+dDrZdHhoRfZqcNZ6
0wolvgNdB6/n+UHdJ6BE+arEJjTUGehnKNBiRC3TDmRXakthvyMkg/bwPWfSQZVxVN0nizpzCeAF
NG97c7O1HiU1VVk1yrXag98Zg9pb9Ow5Q/sZAEnWufRVai/9fBqWuIjDlh56xVvjeyMQI8d6aedX
RWEu5eBCHgy55RXOxZXha1dl8fWBWHvk9erMGjwwRKG0D8xSGxHK5cYlhQ4/imRkq8rdUBQ9VUjL
MC+FM9h4KdLJYwcq9Mjg/L74lUVjjKR3UJPoz16Q+e2gZFi0aeUMjBAo3T0kLRHYTfDPh18u/UWc
ja3cYjMJLEVoK4HvdLJeccgYRdIj9szhea2MVR2SZ5FUb7v9quuSblAOW2LpW0uNHFvGIhC0SCHC
v9Hudk55q1mI8Gxm89TOLhD/1sGd9OdQZpo78OTlYjOPVfdu/no9yNCga7qaKsPUsJAlUuoftKB5
mp54GNkSplQCSMwxxZgnuPBPEkPv8nXoIpQQK/FeYy7fww18XQlSU2tZUwoVEl9HIBfHJpX0ciWo
eTk8c1szCDcvAPK/zOSCLS5N2VL3CSXQ8K3y3o+sNOivg/dN0udaCsPdOAVK41aW7QdQkhFnWIJZ
tZxU1RtnVKtdR8hrzJTpBofqroHedXP5ITuc1E+IQscayN7y04p1uPmzzXpLsg3U1sm66C/9nz3M
UoQuFaa7tSh93+vusIaThIZq4bc2lnp3o2Sg455XiXRxc3TeIbTz10HqlYMjnQtZLh9D+p50YgZd
Tm5Ta5ROEvlIWAn0N0XONWro6K5C79tZRnQNqHgm9iEuvtToKedPNoi/Mue6P0bEp+bVy+L1id3U
u2vWDiPBwjswHjgPwiMRQeRVhxfx2nRYV6UYdV9VZhu0D3G2AeP1+08hhFZRqWPhUywGmBdzgqqE
P3a/UMMcpakKO75PAJnvSwRUOdJNd3mjEUmS75lYZUwYrr1Bag3BTq0bM1fR84x8lfDvDsFaThHK
Srp1WQzk0ezBJR6HoO3/ZLi/FoH6WeNYxGnUYPMLq7qF4MHKsvOe4afKX30K+Z+2l/m/RNhqXoii
kPcguagvVt+Fiaxjl4gcudNZVl4AmZxUp358WqTVIqeFwhvvC2sP/ehDP0grd2/hJw9DvWBgbqML
dNZdhat4+oxCFCmepbUGfbf4sFjamUL3xSDOOScbTC5sLfCAUTN7mMJs+Caqc9IimXBGIAO23GwS
ONKkYQTOoHcZ9VZFi7gFBA7tbPQTzIVccpuZO+alKk1sCxe0IXHQGF9cmtlUo9Pky8r2aRY/o3Vz
qN3ye1ZFL4ZwBU6gvJXtLylsJ5fD+BJ9S6QHApCde1QLDLe3kD075CRtvW5LBVPc/+K6z2UqfylN
CLXJ7hSy2EV6VrglWX/aH1h/Sr24yo73HofxfnKn1jtBEILLueXuJIzmet39hFXAXzAPQSC3FFFl
EdpFcE/M4uVfIn6tk3/bSQXN/RXNwp1s1Dk1ryzrRrAbnNzKHCsJaeiQq2jFAQGuMY1psGSP04o/
4NagEAIjuDmc1Lq9TZQ5/s/KtkmMNrh3RvxnH0Qfot7nLSaLFzy7ZkhIDwd7Z3i6IfEjds3QlaAS
r4Dxwhow2sxpneEk2tKOS2sr+7MDsFhg+oICmWWTxQb8hNlwMPs7v49+fJJoUK9RwVeiwm/uwWqn
XYVlyhDdsJBx2+iJLl7WK2Vj51Wpl7alE+yamI9IxPi0gmlpBBtjRMWjH47/yRPvRdnWUKCPEDMU
QHslvxGlA0StZo8e0zbn/nX+18G98iaWymqctmQAPcqUBKyiRAx/JmrWarEOMEWf2ll5YxYufihr
9ufZG3XvuR9PbqVXgBZlGoEsSfR4hNVsP0lFtwmp+nNj/7DuNbtEjXcb/8zSGqBGt7yh7/k26CbO
m2WjdwGul1Oo5v3khOZNFeakGB+w5F2/dDS0IRR9gE6NH1hjRlZmRK2vZBkgsVUWircDFCFvOjJe
Uj6qwYf/QNYBW0wyeqbSbdr46ZyVM5fOGmo/UQnwjLTnnV056ffq0/9q9c+ZlktQmLLdq9uk3D02
lj/45ER/8ngVzKqVgQN6o+9DvuinFqAMP9x90jL+5KdNs4g457g0K81fr19MgGTy2HdMMUbzEBiG
IPCRZ5/RfH6E8oScAeMRxmEza0kmq4to0ZEds48oLMB51NW+2j39nYINAFtueKzO3HpdaIwc3ZWW
OEdFhmqOgpyuAWaLx8QD8p/YHOuTQWqOcv8VK1wh6oINxu5cELTPHek++fXjYT+PH52KOmGGJaBU
wKHf5K1ZwXTY/JkoVRVOuKfun7nM0MXs0No2qNboLAQAV8ENQf2S1OJ49842v9N/BM4gLfDZnv12
NXmNwd2CymD22kPrwMFPBESOtl7gVTb4cVPLdju87KfPRuAuHwT93LcD5juw1XTDVXkjSfhLP/rS
UXYcBNH/iuxV7z40U8r9CA6ijAHRwWnwwpJ0oGqyg/HMNhetJwjz0/S3VjVur+zuG7DQgteX40az
TEGY7WwnQ2uCB20fTSETdex1PYLZ0+2pKwliT8tDaTfHo8sTzOkDRxWZKkqtPJMNkKn45dotwKxA
U3NIlfudeQhZeDAZS+Si/5FRVpwiVZVu32Oy6lUXluoJDeRO8k5RhQSi2I3Hjh2zv96QkyziEbnj
xCcNZrKdYaxa24WNAgaRc/fV5yL8G5Sc6ogkjQTB6m0yGEqEgXnVYA6f+eWkiHMg5/F8ub9WI38T
qyg3dFEYf2SHFyqHu3H677X1fkfQYp92JS6DX3ITcfT97yR1QCuxsSONUC4tjPzzz53CF9p8moM7
crano6Cos5zwAkCk8fh8Zrb/5n4TFwl0PmkiiG1s6WD6ta2mEeFXENYUXQsvjh4+S4zYVPAucEPI
ftNwLQ5KffwsG9SGlF2wvuSIXYvumB4St7IGPs9+8YaWqaHW8NvuxFekt1YLdrdij0mCHEIVTM8a
v9kckLkHE1zvboPcabWByMrh7R/vTRRX8MjC/pTJW21gii2CaHwZhTSh0pNQJBp1SV+9a3OH8nt9
XVFptpkwHta/NsxsqpQDHNmxYkx/NxaALPYfyr/7U1D/j6holv0pzVPpwq82GLFXyndJzuUFyIzd
6Jqo5BaqtE3LDqDicfmtB2VdO3OTxgrLwkGQs832COkGFXGMOSxa9G3RMwmICfvQ23F+P4hn1r7a
CKhyIsphV5CuJxEhwzW6Lt+ReDxYBdJvkv6ShK4fMBDoZ8m8EL0iFjnqHjRgPxYPoJZb2LMnG+8K
Eex2Jbx3FoNsgoC6QTJ6LLpHquB06NiGVckf6WWFW+Tr0YwNkB48R0Q2/BR/Dfu0IYOvUr+uopFZ
4mtdNOl5dB1vXBfqkdVFvBJZM5fLCYZoXSq37fKq80FEjvwpSnhJ+3WpCPmDP2gQpAJJwqzQAwOc
EEjyCpB9zkcLDB6r+xGMIeImJk/kbUhowi+g3N+VPpk2CkBPWdWc/CX78HX0oUhOf9jSfx0O38gY
u9JYExwq6Qx5FWbcYQgn6TQx0F2IG7UpBrtNsFUcQaxTBHfOlypPMFFtUDTf49MWUTXJKrTbbkT4
tx4ux4veoCJ0xGZxdcqoWW2DeG2Wk/cn5vuxazzD65QRb7b03ZCkNDIzHu9thmNgu6JjvYT7bwQU
wcC0FsMLgKzR36GWHOegcKL4XAfzkooD2iYKAU138UII+KAPzcJtqgYm7yQlVidl1k/68GQUap3f
Ba6rB1KO/JjPzpVDj318Y3qOTdX6tXjsDZiJy/Wi25q4KMQ9uXo7z/h42l9eKgqg8k0eLMkgZZH8
JcdAg2bpl57mod4Tb/Fa5HjuA7DAehwJlcwOz2z4qMwMWRAUUnMMwFDXUSeYZu/fp4YQkaiOSIsW
XGQOVstKr0rnZgDAzgUPpUjQp3O2DBjdpTsHwG/VmR8FmXyYZ8qHIDyFwcDvYPJrE3xI+9HukIJA
93Org9hQ8Lqql0R2vulHZGu4dsxQMWMrlmpFs/ye8J0Tkcdf1sG8O93rtoeWkgx2roKwSVTTZfE9
XBy2BeBNIZ0/4vG36YHWYaJ6gmj30XLRlYQnQ/CvjPpLUxyE80Y+ppLsvNMOzLL23okRyU3PNHUI
870CAG8Be6Sd/tGQLO5AfKzkq/N2JLCRWMKXuykWdER7Tcmah31KOeKAZFVn53O1t5RDrJZBCTk0
SRQsLZS9KDsaX064h8EDLRMv6UUkjou9Z7LuZiDEoProwC21F8RdiqHzZsoMpOx4gU2TfSfItDae
7sSnHMsQUkbvyqz5TYzwGTWQDflCPMe0qSw3wdWfUHndbV1hHbRWmgzo3Q7eAStR1SNN4GGJSB4b
bJc6ep9b6AQSfHiq3xoLImopR8OfZ7smneo8YMzWcxxpkaCLvyraWm3iMbUvqr384YSmufiV9ZuM
geElkPUZ5WaB1FrpME0IpPooCbccWMtT6RZ7FB+8kDB/CQyPTJxIdRFM5Nv56B4fvJIWERVZYhzA
02eok5PNc4w+IvTk5KbJVKnFQfiwhrTYWu0AHkbqZHQFcBgkoXD6B0ojSpCUYMUV0pnBHXm50Wbt
yLrqP72P/5aRWpjdUy8yjXjhZPWxAVfnMd+aN9woafwqqJfVvply8fH5lQwA6y3H0UtQSFoglSXp
KIkizxYaOorE5CDZEzZvPdXhbyTQZ5uqxkHZk6jDE2anYpcUtrYQATziw0h0nf+e5ZkHBPmhzd4V
PtqWSKf9ItYMHGyNHoC63VmT9PaWxSumITOjTqPXIfdl0gZyeGMtwX1Ey8q+y5fztLNHV0o1qLFg
LfVEUcqIGAzWJIaAyH9dJuEI6gTvpaPjzhFfkx/X7emVh+C9enAGN2RZp36MYdz9S/+h3wFLtpED
aYGSy9BumjrtrA4eeuzWpZWX7BBX3epHLa9XzLHWmlr+EVIlQpChk6nm2mAV3wVTX6dpF7+sSol/
9zhasGkOrcqv/iPAnlp5E6A8Lm05K26fNcsLUox+fP/4GXcEP4knjU0aRJc5JfXwE/T0h7aKgozd
hGjCCXQ/86REq80gasFf+k8SYGosLBa0lBK7oHfqdCfPSGD1vmb/of9exCw25vAxcW9Z4iTFdRFG
1MSaOYv/rjFN9wMlzg4SNzfEZMm2XHekTiImx6+9J6vkVeGoPfxlbMoPoI1ExxbwPgA8Rsr/phI/
+vQBmHV7n78oAEFwDo7fWEGHzQjkBcTosGqWuxwiYILcXEKSDcipqK8NUhNgn/vwgMcIzbMj46yp
ioMYrpIpHNBc/o81namdb1+m2EwQ7xjiv4XwYu69tHMgZ8Uxtlva/If7Sh93/n6aQ42YhTnI3SNF
leGD2r9B13rPe94GmPlLHhT/Q1pt9YZfMJ78IZI7IuP/JXSycWlMnBUTCInMQ2b0pBZGT44GFZcw
VEKCDyZGH24UyelQjS2ZWh62SU1L091V22NC5DLOenwuJjIywF45vXEiZGR5e01vHao5wUHYq1A+
FeTWIJhNIe1//sGlFHXD5G4B1f+ywQ9TpjsLdY6DS97IHELIkhSWZH7qYtSGELLmjLn+FO3XLC8W
Ns5kMF4X7fHedw9n7qgMS7IOEcDtnk7yx5e1RIGDQTXeMUoZO+ncqWHf9pMprBbae4fpi6s2RPs/
TnOPGx591bhZwVNK3k4gIgFBbIjDAegXMGShFAvQNsECYxZa9mxTVeXvyuqLgNBRX0z/LhQNO2FL
OqOGDJPxsFhs7P9eCexKBY/u2WhJ8dsJ0e8WYCyT94laP6kDugK1WvU/SL+/ezao66u935Q+yh2f
3j3n1qaLmUomLzZ35i2W+n2d8LA8hH5MvNdvjxliLTCU5qmIp9sRu3k8LOLXnAzuscqRYagxuPIn
PvsCXlKS5sfBvGC2qeJmdAcohoA71GilF2KWK8EvrrNhzK1V/A7H3KbIrbDmzyAfixC6527NaRv8
YorTyGJeBHXjKxr8O3o1cBs5eyq9b4A1oL8Quc+kjLo2ONFIY9XvDHLgjUrBwWOtj8W0XlSTtenW
fcR+YAqqqOEMPNC7T+cBzLRwkE4dV5SLhkwZtU+rxNLe9I3HJwGmIqd1N6TWirycqM7DA6+kn61v
z2/N/mouM4jIMiP+qgofZHLcINlxX+1iqYfJg2M62IVdqEXbu1EZ/c0WcBwKa6K6NoUWFPJ+qCsc
oBWhtDE4WAyiRw3E4XwxBektBemmAgYwVFZLCeWwOq3x6cX39i5aAkcQBLjAzaIRGoINF+Ssx9iP
Ji5cbRFo25Qsim6Td09ihcUjeOWxuACsysofiYYBCexEsIbPHCE5S17wWk5zMwt13o5yI5ZOBX1x
TWHXq8QpOyNv6qloMH66U/H0r1xFzcyIkrJk4EYz7u2fQ9BaEcRhINyQMO817+6bljsYSSFas77E
m+DHrxTtzejpGPYCFjl7xtlny7r27sfjvSesFyloADCtMVKBbvDv65SOYHAnz2HDk8BNojNEHNsn
JgGA5LPEuk0PyKCAVC7+M2TQprvdd1zzdsrShmf/p9fSuve7fe6HdLZrPPMOcfGW2Oj/KR/QfeNx
1W24JFDtFFyjeZkRUBZhWT5UPsi2HDz37Dy5hvvUdmiSIC3teBZg+L2tj1TEjzix1JXXxlT2Qz0O
j3teph7Wy86nscKsCfVP5x2SeP31FhOIhgLbDFym+2PLTUK2OsXlguFlWoNcOGkxD46AdtNR5RSY
lBXhDds6TLLJZcKfThntTyNe3DgTRmAWbUbO4Akmk+iVTIYxngIEPuvWd0Z9HiYqDFiXseMIgWPc
TCJ7xseg1NjrBz5tG6M/8uncW1yFGb8SuUvyv+DM4ESuyQszMs3q5JcnE7BoJWNnVtGW+KWB9BjT
c0KxHGY9cK00cl1SQmx2kkQ9//CNdyjRg+AmNYb4IheA1R0iHN3IJlhfNVo6UtodgVHGfgVd41IE
RABsL+yK8B3kcMegZ+hfmsx78buqlFlZo0i/dFh4gsH2t1NTnGjzm6yrRy5cg0J2VlXg7XNowAj/
TBmy5S6dCcA9P1XrfvEDEanJmbjRa39KRqW/G+wTb72DKVLTntwKbL6bZQXE4Zf/g8hUbAW3WEV/
EHTzKY4Ji6rVlPr1EPhLD6tZME5p30B059gkh5XPGKFGcJyWivUn0olmrFIzz/0/FoYMdsPetgSM
CfAXJinh25HPupv3NdfLECWqqaE1ZKNhf9ZmOAfN7SyV1Een6LoX4BRntmzeJQrShl4V1KlZ0bCJ
U7NMnOnpNa3j++4QS1oaayla560cZMTr0feaERDiFEb9cf3lGH7jJ5UkKXRJalC93TMmh1MWJ/yv
84Lnn+l5D67+DVrSDo29W51gtscS1AF3cKtNByUZo0t9e3zoBNpl899DjixN3Q3+eoMYi6qTrQz8
RE/JdQCunY+343ZRq3qKkaQGvIRFT4325ynuDWIFuBjIkMPCj+PUzi02PlN1LNbu65QHOa/TcCwA
zo0nUI2bZ06jvPMdoHoFIyXGmCji5eNWIQd6DAcjw3W0ccxixoraLBF+PSFhtzlCMHJK2KwF7Y4Q
a0rtzauwemh6VpyacqlTE9EcVzjuXJKh4bSmegA+Q7It3v+7hLL38BfBceYSAFM1wqHReJ2R7RfO
cvWZTabQ7ezNaRi2C4xi343JUJYPhr9FRJwbZbEV9gP84Nu48W3A0RqcjzT6f6hCXGgZIerUEW1p
+CTi7E+kiefBK7JgPJkd/f9eQuq5rL3eL/pB6Vfz2r245h6RWXecMi3WpK9t64na4sA8TGoqaabr
xsj3zYn2L6v6yuaXSpYs9qYxhyRzmmcRXw9O9YWX9GdGZiL2lq8AI4YBEiY2NI7ZaF/nyKa8akfv
lb/TCjg60RSSpDgc8KIWh//P7sQXbCRFr13ecD9nR1x4z5wZJXamUKUXD5qXh8D03rLoTwlrcZa7
jJsYODe64PG03TRay4EkS+WLUMIl8A+5jtfzuz4EYob++78KXJfk3OEhSdakslkvGvDai8rvcniA
klRl2huvoT60PXYGcqF0ZONCrIt5ZUSkyfayJDU5ZVNAQuVTsi5o/OpUOfiiyAUKerC5ZGZGNGPn
ga97LZh0s4SBtCa4ZR8epPSiUbQNppyhj27KR2uXFuF9vuxdFRBeDqlVR3pjXCVouuCQsLixi+hG
YksJ/0U9npdDDZ4jM3TSgxzxbjm1xAPDUVhqm0ZQu0MeUKk4ybsd5yYUaSTU3bIUhxkacUAN71Wn
CeA55bKGlAS/RDtzgJifYcNhRvEoHEyfIKeKGVntV9CGJDaElPpOFNGy/K/oYsy7gICcqqz8B5wq
Byh6k1SDP2Fp1WEj6Ta107vE5SNxz3qY1Kxk5394v0XEXEHIDcHO2/USO52NjISX2pwm2zWlzAhb
vE+HZytUugVUG62TypB+iWJh9Y93gdPvAFxLUVKIxRlPI4/t3osFRNV3lpOsj52bugrmoioAsTNL
eCg30BHYrzd1EkZQmMOGJGumP5gtO+bRSHb4s7RcS3/2JMlvwHRw88Ov1i29f1KSVhEkgwU+ox8e
/iySe0dclUMqNVnPtWF4zI/cLprf3dwnSjamgD8DLr0oIrqIQTnq9Gv2WGUrkg2IYDLc+gkppQ0O
ZlOKh4lFHwHeDZrC0hd6aR/REVEh/BIR+ngUNyPBgbd5QKqzWtsR2jirLeqtHcTRhnj3JGNmwDrv
ywxak5oZ4qrVj1lpWfArZDbxAlZwR3/Y20jQmJACoKkQymg2O/DX91+LlUR4EgFvTMQFSuFSuKrf
FDl+F1ApqvkFaiv6KH0NSACF5Y6Xf7G6wMDU30v9yxrFJ07ituPDp+TVc0mGR9mI24HpZzjSXVh/
votAVkDoKASqNIbEol5DyE8k6vuEOB4B2Ggs8mJ534Gw5YdiLM4fDyYPHxbA570fI5KlxwEAelZf
w5AFV788m6GDTe5AfSNfuDVxZuzVgrbPBFDF68eJsyk3ne7BKWbQMtyOXAZhu9lt/+gPtcy6ww9x
QM+yuipIJ8H7rCaFv8RNBbIVrR+bhn/x/7mOugwPO0nTEN2IxePJOEzQjwp+TaRhcv/x2Ku5zXXa
pQKZy1VltH03welqzNmIroAGqViLCr6cuUlkfhv8K86ekrqz+ZAjbGUjuGbYdCIg7y9ovZCeKa9j
YuWkKHNitXlQQ2Q4N83TApYqIiYkEuwmZQ9VieaLy31y6fo4OMyNG5iqiZ3M0sV/xVTGPj9hX4Q8
yGmPuOl7sWeGrKrMA6DqwHCxGe84RM+xsrLZdehKYtfVTaY1lSBSGLa0Kg/7Om75Gpj7XiOmY0nE
ROyd09zRqmS5JGV/rNqmwHVumuvKR9BYxnUfj8w7NsE5KRZmsYxIZWARjnDns31hU55EIDDV8/wo
ORCYQZoZO6JRGV/20z5RZ1zSKVhdAMqvXZ9T4etRXuwdPozJWcA2piP0la60GfsrXHaJr5ACELVD
E3eeItLvX2vXC6zPNu4tpXExlMcsBvKlYZAX7cM6Lu4sAzI4K2EaV+rA2ozeLjiBZvy53wJ+AMoB
MKMF28E0if5/Zvwax5M2EE7IwOoyNpPT4qTmgN5UVzuVroJGbwk6LELwVDmTTk1LnLc7Z9JVgFOV
pxvGWBcvEJxkiwl4RyBk1H7MooOJn5P6O+Qlvj3wUPu38TAUQxsMVlVyD5jWDQ/uvD+gKQYlXNU6
AC8iYCrgs4yUZR4L2xt0roDCylZ1OtimBL296WNE7jz9r/cXunm7Y5ljy2L9FAdBEEjaOybn5EKb
x8OipEryLXK9INHNmYyxamqbuTHgKgfHTgvwnXO6yW0/3btg4kRPKFGnqQvPWKz6X0+8ZIs/jldI
1GZfYZBCjr83W9hEUEEEh4MaQ0rpaKxU61VrhJM6NqazQB86HO/ApRP8aRfLurLTAX2Jt1zC6k5q
fPN79GRp9qjukxK/AavmSAkVlHxYBPZkkK9zz+zZRC7AacSEg1xe9hOAQGuZRWCwCFcZ0+jN5BfK
pK1I3GxPL3d9LnwbljjMeAS1WDZ9F6xvVh5J4scE+rmVnU+dwKwZJOMjRYryBRMqvEgs4L4JTgR5
zuGsf39oyIiTNk4sz4/dHmOrGT3O0DPW/lsZlgu3p7nKCvcU1/AvEDXLfZ5/KjzO2Bn2pZFa6HUn
w00hMZY7zNxR9ue5EF+8vU2X61RNFiVkgFYFGJjoeElGUgtRFmP+Pzr81tk6Aws69z6nGq2S1Wwm
57ockc1g1WaJuPAzX14weara++/425Xr19HzCMNJa+ioL/lgtxtGGb08LPf2NRG5qLP7iOxOeHei
GhEzdaOpuh95kEnPPk2fgA3MQfp5+1ASqY9idOza/SzVygd5uYcV8SzHktyDHUuz+564xSJHUYhd
Unx53XgdENdH6q/UtdSQ+KkLKfPQ4ro6fa8IpXtriK5vjrU7TbcT7Be6a4vXU9HYaC9z9cUbA3Ww
hSUTIyLjtMyw7iqOoSeGCg2cfDf4d0hHL9T+BHSzJxBA+UdMAePt+gSJKyFyG8mA6/ovsD2U5BD9
Md879hqzNq0VFjUaI5kPM63/SrKZfrKTPvMV59y7GSLEFoQoyrkwgNuD+O9fAKw0KtIs3swTnVyx
FD+rtHMiZpA9ligr80xAf0+/eCCKPl2nu54U/md4pibxkkinK+TEITcuZ7AHCmaAxxMFuYwYWTCY
xePLR4EuQ4jriiWZ5kEECGIyCJRtLM5S2NWmR9JvS9BDz/fiN0KDMwC+D0E2CgBJypDMjjQelq/K
9lXr5zVeser6cCiRwkVrhSrRP7ggUdPhS22QV4Wy1zNnWWU+XYWwTwVrbCVNEetumHnJEqMB84IL
JPh0u4lQosEfEwKjNl8e9FcZsO2PXe0eGQKZjCAOTCONThhgPMJXDlWiWR7jzHUqVUDBHEcwvZXJ
kKVWY3MRnaHg8axDq5lCzSS/HUzkGqnMIMuiL3y8lVKrHvOltavGFewqXrQvWZMvc4WSDVPqpKSV
ZXYGyInzgm0nk3N6HbNqhpPBvvXBPB5jUa41ksHqzjuehjzExhMHh3oL+/+3Ll35h3kezUYDtQEf
y3Pjeiin49K3M+gBqfjnKbukWsrNYKuLfzZLNZduVsSaGW9Vur7V6HfqTqN0STwNWSEno36uINFp
dTcF7iurEmq1acoeIWL7B7H/0LzIz9gkglStYtYeyOVVobShSw4oX3Js8+8n6C3xanTxuNQ/DeoL
Xelc9v7vaMP+E3SiXJaO4B5s5/9ZDzPFTqh+RO1KcAQPDbX9hsgkDtawhXr/VrJG7Kk3AWaL6vD7
iiFcM5WdKBhLBQEH3+QW1OahH/IQ8mKBiEMjn2hDOmLTUpV4jQcd+zvnLpXQcTJ9NGtZpGpAt8OR
kgkQFeGxPb8FZ5HeZbgJIr0p0RECxFO/uDEXjTRFw8ZIY0xttlVYvMPhgrPtnp3x2azCD+7A7Wmj
TGIMzZEKOKOWtwsgW/aaRrl3rzYq/4nyJJ0XIK2NTwY5y0UwEBA6qo3hq2GCrG9GZvWoj7tPERda
3KLpDecuadyV8qxmo4BdPbLYuYZwheJMom3wrSVvDShn/fA4ATMjrEUd0uJBU+elDjjhX0uaxxC6
fHkmIQknvCJ30MiTw21ymjG56Vc5PgkC0YPs/tV1rGHadnMhmIdVWbBmc2KW7/pfoZDwlGrdSKbU
nbEyuwhETEBxDaSYCOyMVMVOlkHpdy9/KvvZRCzRQoq1hgIQ+yjkCHcbhGD2HcslS/jrgUtGoRms
e6Z3dfcmEKbeYVhxgZrTGHLMf1mglH9whjBeqeq1AvV52XpUQuZ1gSzmvErWRRqJCKl3MyHi0Yhd
3BwPm7nXYjVJCGP2hGUorVYqQGcoxbbBmW8Y1ItT+TFf22gIIA6XaQTIAdOZtjVEaRW+TCJXLrj/
k9cBcxhgh2M6l62z2SDiCjdkxV0Ouhf54tCiH/kyRYE0N85D0E48ASXp6mh32GdPfPKVGQyN8ioA
QUgMJ/i+Jqa5znNu49lFRMn9c4PabmO4l1qtkqmJ9RlwLDyjL+syTHZ92ehUQZeGskGrl/rDolqY
P5q/dN3rULkkW4lhNkO8xd6sHUYzlJpKe359w/nkioT8b35pkcT7JtS319sOKz/FJepRzWuTTjvb
dCNd/Xxl/DW6wpiPnForW1SWdYFp6G0WMt1GFbCeteKwXpFF3fm06diHUSg9VF+L5mriASpFd5BT
4s8WOX5ko9N9oyoHSxRm5AAAJojvenx0Ce7Ki7qk81x+g0VN2Nl9V6C538CwsZAUdSp1+K2B8/m/
WzQOXYAmsm/BlcVeiYpkvoUhDnJGLPtyxwY07ACijgkoUABZ+YleD8U6aCiVYSCTS5r5MjlJaMUf
szK/vMaAppp4lRXYKfD4ndQD/+QGo6WbgoOB1vn41pOi9cr2RYCjIocMBdosshI4FFsuDOoZD4R0
PXyS8oN433UVRmOHht1r7gjnNOWmyxxcIfpBWl2XOPRBSWN6sMk90EIrAWwgHVzEohZhpFv06JF6
8Ysl69eg/AvDZTceE+mW7huX307H8H2EKK8YG8AOI6rT1/GkhqkrjrOUA0JbjfokJlxMmbhApxXN
GAneJOMTyOxp+UcGdz8SW2k2QzF3S3Pymartt4jTRZxuR4ShmHzwLpKguohustC5weqZu+sTiTE0
mDRMvkkDr2LyFkn3iDZf2blaKm82ISPs9xiiKp/hvPQgTxTUZ5YWr1fyd+N0Lhm2JkUJ5APwbFiF
9sJHptg6Uq3lxqeHpDaMg8T42K53jEWRD3D0yZ5RLhQYDXve/KeHHHw8FlAXiMfNOwwcepeGrOof
dg33gS5l63Sp2dylfrVsKnmapa58YEkTzwRqxdxSm8XopuU7qNMzqPIbY+aDIESWBtxxp1G1GWsz
I7sW52ewZv3MG/hX7Kabf83/dLqY5+/0YOGXEGGDS3Dp2r1gvHquujSS08tF1Ug3ydCgmilVD0xS
DVY/PYFnGZXDOHbq964Fi4NlHSt2ZclbUiLxuv1Bz3Q7WeNWzmUQjRzT1mKHM1KWF2r/qvMH1RlF
80kwfifExLZVt88rSdoZWFqAh5OwEPNGIZcNvs1N107AJPhR6ky/iOJy7Hh3twJNJMRuRjEr11VT
yGyhWQDUcxxk0bWY5ZKHtggWdtEvhluOnXgLUKtNSZmDtfMdNkNwGTDtX0NDJH3CTim/aqK7AKgU
QCdBYF95TEYi356vnQmNM4I0kvk+vgJbXN+OZT9OGc2YOzYl9n5pD7hh2k8CrlmuAmReSyULU6pa
nvPq7FfTzJ1QybA0UgmPMzHWaq+tMs+TBXM2mEbkQsX7gqlVNqxewF5jOUmNX9CBrebkpUdBDP8e
bsNhWI8zLYJTjhMOT9muiff+XBf6/gWF7ekl1v5NnFzOWlV96KgvsqZgmLYCpq55izDVcCGjVMZ3
SgUBlBepgUi3MY/p9d4lOVbHCWcUih0rhU2tyZzzBtT6puMz5GFVO9CodEOWIoncKrSjHeguZh3u
2241JsKVMrGPwl8jsn2iPXnaoqW+TIH900G/9WwrqH478Y92bbzvMKr6n+VTbL2cS4h+t846qMWk
04y3PQUL4dkqu5oj1aB1Vosml+uv3m5QosFiPfWIo+sL8xVFaQ+bMmf+HIGYp2cyyr2K6cB4Pzhr
kWiQL4G9cB+Rnf3qdnVYnkKRURzo9nrVKPsNI+EOHNcbLez8EtkFlKoRnt3FCxuxV2EKgmC8h5Bm
ZBzup4K3Vj90/HyH+UozI7ClBV4Fr1CzZ4HvBdsWHipTxGKMvg2NxyCHGO/lKbCdAUfLdV1lglvE
vBzgXgZ1J2RzcktbzSBlxain8P4DrMG+mEt9f/YmLgoNdRS9RTIrdYHQe3YZN5DBVlQH4ICTi4cH
CrxsawIjY3GrMU2eYHkc+dTjLysFsXaemby8SvJRYUDoB371osHX4+3soRWQ6YSfZ2P3M8gU4rEA
oiBhlzJon+ptB8jBoRq9N3x+QZ4XpGnmaS9NbjK8IfoSazA3JJas5dVc+VrhQtv009ewoaZ7QWNL
bHU/yYVb7k5qFeAs7735qve1wbjey9mJq2JT6DEF8rlGtv1WGwtyOlaigcCcD/Dn5lfcHq+eEDxB
knnlAmPRRqFqC20Cy+msLP74z84Z4gOFKNC/AOJrIMIZkckfvwFGcdDf9O5aaLd+/ziUoB8qbsfE
qskQUSpV+9mS9ra+eisUJ6q+Nd/HuzcyUFYk7ij/+qcctVN2Q73j8/u8RBJDlOfWqEw6bVJjLs+a
geZhsrZWhz/CUVUZC58iWiR18i3ROM1y36Z9JL7UO3M3tpUJi4sxU+SNWyB4T4xLVFhFusx59qA1
3NCsD3SwlDgrxHhWyDDU1USFgoiYB+VYr8OUfU/mqfNf95iu0Q64Z9q44iUIYbkcz4DuThsW3KTM
kT5ehBXgyoGdcXo7zbzc29Fc4aBfuqRMPx8NQ/tLDDxvANenFT7cIRLU5/kCGuNascRSpGwErwY1
Q62cocb1ihgdGgaE6wiF/5HFlDRnveLbeMVmNOgK3QsaoIehpXMsKeLw87ll77B4Zo2fntQTKhqi
0gVr6qWniWFEBmWPB9Vwu0NvB3eFD0zZuutih0213a3zdgz+AksY74r0YQJwmOhj5o0XxtAZ038p
MAIHYTHd2nzyol9QxNGYbqE6xRnReHGRsIi1S1cFDwkZiEcE8FkblERtcLpWuFdK85I+EapAjgb1
soS6YQH+3qWMPhglEv7aA6/6T3xYX7aNEd1uLYPh3bxBPfXr4WalHPD/uaeygSlPqXQWG5rxUSxn
M7kanQ9c+c4Jz3Gz7Yx2MnmSp2vwLtkhYNjKdB+eglkWxBURMHO52XZ8sw/foc+IL/W78PheeD1s
UDVZZgN9Pl88r7NhhZGpdVgoDx5IZ5dhNRXwbSzibxNIbrfWKA3572hFwiOGNQisqGJfujQfhDR8
H9hbsGZaeuiwvofsqkNdeQ3W1wy4GvY0DCjQoGLiCnWLioc+PYPCyCQ9wBcif/nHj28mF2z5jDLK
yejhe0KeBbI7mCfGX+b6qljIHHulX1C4XzTS47zxfcfB9GvNeqxezFmUIsm3lhepmFQJvLQOiu/X
pQsw7Pnj2TSdD+Q3y46LCPioi79AzVLjgnKtbs2T/gNWeGxrnFMV0moPHA4GZ2Twu8fDA6NsrtHk
F5aXamVp/qYwdl4oJSbj+55ERQAMsXhsZYDgJAs49tbBzO7Xpg7qU2/Ke95LZSmdEC4c7kBLFwsz
vsKECYBQfxN4U3+yGahKl5aekGsxLS4baZsQXntcbM5ivtlPob+BB6MEMlBXqYw0ngXkw08Yrf8B
A1g+zn9p/640DiF0D++hd73neXbhYAPbK2CAouO3L5h2k+4aIHzwVmbhxh1VFPVvjilaEKZBezEE
H1cAXvYbRbDo2P3aUdn88goaDPYvXcjgcGC+XaPFbRSjJizumoBFF9fN2PimxREpWIHghF6K31bv
ssfaFsK89ULQ32z556uwtX3j8GV8EUe8rY5BLacq3Y+Q5eqm7ZMTVBG3LwdVN8HRChB5qubpaEv6
mE6ou7JmC2FZYF2lelpmxDzMECK3d/H5jVTXwJQI7xBKOjwXQPmcjYFHoAHrmNs4qbD45jre4P8w
kAHHywW5x3pefhimduHB8r+UFUYBjXCN10WkmC8fFlusD8yd7bAjHN4B8sybvrZP9SPwUb8gYyA4
Gn/Tlof4k4/rrzOZwXrcseuZAZ9vwX7yjYm/KrvupWIP/TXzXmwQI95neouppD7RD2lgbFaZ06nQ
kcPrHdauXYX2H2rGeWB0jR/Qw9snHB16xrqqdGyfk1Zxrl6DDjaXU5qbDIvTj8kh0BJvpUp+Hp0G
s/7Ub/rDangnQitlmjV41EcQLdU2LGUd8VZM2yPQtYz0NiJb4usQESxXeeb51yXZWe9VzooT0fBa
rkcH1aanDGOBxSg20ROAAw6NpaQ5Oat6Vaqb5ThFYZHjFE0Wx+RyXwwAhL4zSnFUqd1cUooRRvGG
LijgUIXtEUVvxT/eUvMrOtnnOOjf4L2GEPcqE5K38dsrB38PXKdD2H6DmAFlkCAN+6b/u2O9Oj2A
C4qBI7qGUwFnnXYZXiMGSQ8wbsM2ltB5gD1tKZu2Q+JRZ5IcFBAwt8TcL73XxM1v8xEp+7mbdudy
R37UrCZ+c9EY8AhkdRa1lwJzYeWF8IQla3f5XUEg/yQSRVDZO5CQ6mWVEo4d+1i+jBuQVpM4fRa4
lkfGsWwJB8pPygtVO/+JyBcAuKaUq47dhJcXafukUz0oCX1DHeO1sKRRaT4AFr/4SbY6AQlYxuDA
WEas+vdKMQJAKoVDXpW6MLBtWT6vi31rGIHZc9FHxvraNmP3DFgQ4TOVqo1niZnDmix7/g41B7Z9
aS2TdAL/wzMHRxU/8hQURogINs2vFq76DIl1oTlVKIQq1NiDo5De0XSad0unrjvifm1pmcovHhGW
2JHmhdDYG6Yw1d+YS3CqpF4wKvDiyW/6dLCdRSnEaf/qftj2a+ip6rOsqZoq5NickNqkpz+Y1S9b
giLKcuOjXWeQvzAdxvYdsKoB7gRfRtrV4/Mo4wJpX/5bEHp0AWg5VfxBu17/YispupTJnsjFZKPa
CFwdtTkThp22uycQYSuIt3s0f8IMkCl/BuLi/+bZc6tiMVlohYzzXI+Ki0MotLfcJ5nheILWv1Lb
kBhMTRlUIvNoEs0dVIZ+IbnMwTr8QqSQdbIu5THI0jadGMPsN4pHLbSb5Iboip6dWjv+ydTxOrIT
zXgrFLe3ch59WryvUGsXK45O0+cZp1GB6mosp3boE0cEXru9JPYJzH5se259Uhgdxof/mx0yzCyS
J2wJH+g05fdK1TLAFWARsR6hs+R/iSB3pR20xFx/Gg1zRDyxqxWbDfghnwn0MqVkJNf4wBRhaaBf
dfPeV7B+stxVxvc5SxFtaBXqJwOSFWMXxhUmpWHh1AhOvmlTBgBXEpd1j1T50TPjvomxS48FT9UZ
AiSj/fS701gz0C7q5+bu9lX/Jr0G8ubnoiAEmFdrOKzsRFMyQ30K74+TP/WbVpNbLWwN6Y85KR4I
8FYolYiVN/y56dRpsBxVACWCYD8op0GYFQFnuHgxC9BfqawXun1CwopH27yedygvj2TeGBestrVT
saxdZ+rg1s5CyORakXJDUSY+SazRBHZRXr2/Jyd9gMMpq3LQimQxOEL6p+E+sxHseL3C8bgjKsg6
ghTTA9cihI80kZUxLxbMisEtMl4bgoBSpsmHn2CHZlWG4soEEmwBe/nxYpLnW4m+mfn0Fh43U855
uaPrRBBlF3I3pTjQ6b+rsobDeHdQmc27hd/e9oaYCL3SCtcMfHX1waTfHHtk1CK2RF8VY12HQoxb
DrOuct5JmbsF5x7OttvFe+JwnpiGJZnXzs1yG0jFnrqiETS83PfbPmC/X7SlgUBtwGufWglcEcPd
+gZILnb18BYea+irk4UPks2dYBIMmyUgnI75xtMTrAOjeppa5uSfb6cgZqmRhiZCz5TCZvhqAlGm
98DdsR8X4OaHyL/Eduoqzb+krCmN8yDludi8UhaYa6Z8N6U26UDK1Il+h/e56TmjFwQGW7aiahno
NotRyClzjAmqVkX5QFhBky57AQ3yb4+ejcy8vPvaiz4yk0lCxhzkyWaT8gR5x5Q5VlXADF1sIkKZ
J7mYFJNF23+1tTkUTfmgfSeeMyv79JQL83lSqPw2d0V9qOCSJ7HEfW7F0WpU1IIXbSNNLrywquST
Dhtghoc+Zc7o4RMv9ciIR07qomK7p77QhFzq8mPZtI7cZkeQJRsqICV6a9/CLUnlSjQ1EBvUix8O
01eCgSaSEHDXv5+5S7G/0t10ZH+yAWyo53sDqPTa1CKWByi2c5Ns5WVBU2Qi1OZ7gCGLrdJmLDfY
3Gy07Qq9PoIXnZigqxzVFifBfhcDHXpHT8qAfVOXYA7gsWQlPngqQvhGt1FrLDvdnbSR1KkeFSgi
Utk6M6Gs4zOgWHQ9ssx0xu1/rPiNys/PYksr44uXTeYyl8yBmlcmwi3ZmkyhENZqQjoBGK9zDDcu
/ZBG55gsqt7Ehe124/QZp2fgqvBT1tii1NDwrHYE4RW4ztV8bYGFQJVUC50oCFfJE909rCHVGmXQ
g23Xg9E2JRq02mg7LViRxHPFDgWCQYZcMbCppcAg67drVQYBicsZgMcRNgg5rqBY1sgZaAMm5voZ
4HqFM2UN7iLjM9AzcSmXsYG7HaA3PW8tlVZYRqZmzvEfwZ9+FsqLeH6efa/HKkVWNNMJq8gPLc8J
g3sGCesyzxuAzP4zye84w6cRz4MFV2DJpVxnIfeIpTEwqTgVDK0dt5LAHhLdZPSUozgteV6fpmc/
LILd0Cg6PqKq1zNvqNoequPnigRZzhC5RfJ+1XaEgQiTWOI7uSpGfPVkviJDXAg+si8qNl1FHzvY
5dtz5gM1a9j9IRKSeWgRy5jWUrs0PzD+J0Ngw0Cz3xeHrLDFipyVuEOpnPlora1h8bOlV8ElzUP7
4zQaDxcOWMqEkh2HjfCBi8Hmz5LoBpdWWhPAlrQV8msg0a19ttfmST5gcP9q0FE2CsX6VUCueMRF
N6IKDlYRyXeKsYDn0o0qGoHoHgiiWYdvZ5vS4NMoPqmGb5D0xuz08eu0J+j+EErok+tsv7hllXfA
T/oRa+ig3HTIRtLzLJnF+1nhzerU7dRB8hOUgAVNX3t+nXUcHcucro3bXjYE53p5skM1gy+3vLvZ
Iz0fV8DTZ9cf2w8i+OIZ0AP3+9A4ZXyma8gxX4T/PxzGIDzvK33U4cHyv4xIua3G7kPs/T1+8tIX
PPMuuGU/hS8AFMlR4kK4zVSdwgW8dMtOKG42UwZu4DINX7Cb09c4Qf+3mCYw72p/8GXJ1SwoDUBa
yJ8LP6Cq1iNQmS2wdyahoZcvliiIkwtgZ/+FoME3WK6IzZYEh78Q7l7YW+sPhI/FykRvt6d5tnsU
+ZWDBjQvYmpQkpVj4M75t8zVpBiKj8Af3HJIbab++9JZ3lT+dxVGs+bOhQ9t0kXxzBInUu3ipot+
7LBf5xxz/VLPzbBOuC/TfeL/miaEUNkKvlxVtVMtDphgNrjuJuBRPlpcilCxj0Oug1mW2X9HG81N
MsFmjT1pGu1BeoJzjogYOa3Oes/fiphSU0uRO2bDli5slK6iUV923sxUHCUZOAuuF0Ce9RCy9/Wf
9d8gPX1sGN0puO/16kQCcn+Tv8i1SKxxBA1iZ55xtlXpZf9Mo6dFIKgMkucnI8M6qClhkgPDbSxC
lEECQKibVNV6c0AmSvrSUzMBLJFAT625KTwcGmHG7mOAxlrqZdIJh3+iHYp1hfFvtzmrtweUfqFj
RuLWGC5bc6QBhk6me8BwFZPojWOacxiVmU9e9UiMuiWAmLjLWSeDcP1b/bbZu67To7gSAGmD5d8G
SJFaU2hX1wt5gvowjkbaGo2BgfjJGSS5RpcIbMmPkptcHR33VqW5uzkzawLCyr5/VIzDC2HjG3Ue
rppiKhldidnzggZfo3mDhvHDtFNFx/BYB8RjIyjGWJVLQpTp7/cVkmadUHG23Rau3//Ums1CQ/U0
AsL1U651aPpxe73NiSDbLvIHrDsQc4PHA24Kvg9sZvnRTkxJknQ2R/KNkd7V3i+BTqweKGzJ+tem
GMh9Sv54FldT93NpjjgUMNjeitQI8joHvKZckw1jF/u3WGV8plkYOkJZ5dcTR6i2oYC947Qjzz/j
Li8h+6sH/bmfLEvKZLdWun01Xtp+48gJhMmxwb8O3PFhcFs9zQSQqAIYAPCRxrTBI1gOtFpZL3Qv
wg4lP6ly7/gWBNvCJQ/7WnDra9zwi5j8z4xZPyujPdRipl3BJ7RkYw/TURdE6gfzxxUpj1iJjg2e
fJINY/c1U6xYG9Bo5IqKviRXVpC/oRpIzpoS50DBaU8MTMiGo6CJwqS81QJRT0tjgBaxgdaglmF7
Gpwzkf5/rvATBY18TrpL2hK4WKL1CikaGmHLmO3Vp4u2Jl9I7NZRh6t5C4MA2AkgL36545DffkEJ
1Ugsn2fb6Z7mO3Ei17h5Jq4HVwKxQPHWxwRS37pGqvJzgJZ7rBjU4t7Ucr8yybE+IEHSsMEin4f8
cVkUYjRW2Q5ejhkxVBFdzNqoMRSNeVD+c70FXPKB4X6wg4mEMWuROTsn3UOGseg/qtKPsMwP++kJ
BroLChkV0LyGu2jF8MMMsK0m1zUuFg9IplDRmG1oPIy/EAajP5y7j5Q97HLcX3G61eMSlNwlg16G
LzhaHkLf1FB+awASbDCWYHMIqkh3qquQ5WCjvOGN2omeMPP0n8nZJyGfXYiX0oO/A8LVMw3XcNHS
6+VQGWmhT36S+B0u3H2wvlcGPqTMbCQl439RDigL+exSbBYCLjipdE1wEgnmAAHO1/hUyh/haL5k
WVtV5yL4SculObluO5jZULOTfKEgJr8OoUa2M7knunGrifEeIcyeaL9BXKcdCvsQf0KNaSTcz4HI
zAmVARzo750aHH3k1l2aPkt2h8vx7sek1AqXuZyD2pZyzDBuuVE08aAMayTLMjvL57RgJ3aG6tuc
Bu8P8pX9NFeukXhtA4UiTBx/vkABFXUX/X4B2X/6rCtxYzyWzOQB3UBeIK6jH0uQbL2i7hNcM4Jn
XI/NtjXDE7QneptlKRz1g8WtDAwin8rF/UVx5bB6I81yhZ0QcbeOiezCgTwe2GehdXzk2kboA1VE
BUf2T2OYJ8NcS4KUTgt3pV/Dkj1/Vo/gQ11grtsdQXzdvg9x+OGaggVu+u6VrvzFNmcgvrmquIcU
cNSYcpP6IkwGnkw2YE/yfAQG5laEFAqw4j2cwzyK1MG6t8Cw9vDtJuYEK4iUQGGOAo7+qRUdC6ng
khpnVNG2qdWBATWeQjegVaP1z1olrm4wkmtJhyKDeQ/fFTi8FPSwewU1OzT9DC5GUzVOYMDsh6w+
sv3ct2TNn5Sa/0eiNcwkl4fo0dh69N/4F9W7NHtZMiZwi32wuA2KMnulHWSwdcPnf98OzzOdEoDV
3qs057BOd7FRqQh5D3MaIiQYJKxgHk0pZOlRpHQqnHTB4WlGykVXS7OLqBmH6b8YcQr0MsLuhVpA
T8EM2jqo8PMX4GuonMZ0BFIUukx/HFDzlSvshWKfASB8qBdHsNaEwkTVkDN3s2JuMe9EOWrEJarz
Tu9fl5PSvLTa036K0IOWQqK4ZeSK47k+HrekBy1WO/whYFFM/sHHVFPnAj4W4QJZMYUryvPnZLCR
PtbTcFRFEG0IJL0Rkji3Or88c71B12kUknV/LPURVvhvn+v+rjAVlNhwi2Ofj4F2QFGWlfQrZeeQ
8LrnBJgF4NBmH3Lhb1O097GiyZSqce/ynIaKWlALuaQRVdvRS9c1COS2lwAMMG8ZfflZG/fwjrq4
UszEgLRqfr/hGh8zYKJIKXzvk2kpgX+5V2XCEdrB2SBmtbdP8lO6IktpGO8UncB9obr8tcEEPr9m
v56SLBKARe0uUfsXaYOzX+WgOcFpJFn5RTRLfMcfDNf0ebOkoBHTuaUfgL3Clswxs4xPN4YilH6P
6GQIey53K8Dn2KAmqTDIxj0Nfgm5BiHlkoLWXKt7Pt8QWB10NyckcmZ97dcg/Z2gLZxYF9DKC6j5
MSCBZTF1XJk98Fo8HyOYbCWdnkGsp1iAve72R9iHRvDoYlObe2teJpOnuENw27wOVHDa1rmSsqnF
ZEam525+cR4FGW6hJPW+FiEt+2ML0BzHmftVgzUw6W6c0PXk7BsmRykLZVhmVD3IVt8v+JGn/prs
HhDrVJNKm/N3bzi/Mi/iGamVEOwPslUlJ4VtoRASavB/v6gd8fOWO/o8IKCJKMZY0sJxWV38r6XH
LRTxBiGflHttqqAUNne3XXB9WWNm4q0yyszofqZQNd1Na6chX+PobjfxeSVXpxTGk+VjxBJPi/UH
9Q8IFmSWGn6XhRGfCUxBOLhuAat6/QneooKoa9xmpyj7nRtUGnYIstFcyrRUdyRkj+yBUe8+Zp+X
1lqoFm89hyodsKKP4cNjRpUQVTBTN6M2Al2olxdjxc9vBg/qZ6q7eY/mKYAnwiecB9iYD45sIV5S
tYdSRIa6y1Kg+YzlDQ+giDqKA++/dlH7rPkZkKaGnfqreIs5sSuqFvzZAT1n0wXS2j/KhniaKACT
tX54jAtORm5BXgcsHWKRh1Y4WAAWltB4rillaMwIuJQ0Cjpts746CcJaaiLqirh6MK6UNGtoU/VT
9wCv9XXoPVYaqGNBkmprq4RNg5g3EO9lAc92YFYmV0W6CiI4hAF3s0pf8nSL7nyOdd6lgt9r+P+S
K9RkJx207ynqUQmkzQ5osAnufn5KQ8Jhj0mNnJRU6KHykmQf7Ko5eqM0f14RNwiWQEeLrroO1oh8
LuOev3dxx1Te0I++dGetqNxrcv4+RM29pVKEpyz7CJpyGZcqspaLDv4QU2ljIcUFJTHNvfZTfFt9
5L/tNn5cig6HDFG2rZlzoiVi1OZQec89tmDGOHNWrL7JRfH9O35gsFATGBNDwwhrSWnTS6rVZG07
bxbG+iIs4B9yqGcGeG79lVdXIo3fKO/RGTsKLxSDF2oQ911QFYculMLToEZb6c5Xft7+iWYd3ToO
u7R9ipMkbHCJaR6vH/aMv9qX6JNhqLCqdMFwVC00lC0vg5AqqO+yXw0kqtwCqfX0esWwoj35Ocv0
7EPjmTNqDY/fr9GaneLKyistwhSDFGNb0GEQdeVdV+crgbM057z0jERNE7eiTUJCTZ3GbzjevYXL
MdtMWWp93SYsshihytj4X1pJk3+luQVw62zx4GqDiKc35kFL5/hMPMtqV8+k7L2nqE2B2VQrpUaU
I+rAljGiwToP2o/cpHnLxw8hJ+OshY6UGCGdiXHQ6Due0SjzKuP1mXuBMRXdXERrV11z5ay0IF0d
deqBNFRHuBFYYOLo1FwwdA+YqTzQT0XIKMCTvhaw0RhDkbEM3iCJOtao2wmvyl1mNQFysK0B/n47
O/4o5dJyLX+a3No4gbriIO1Ug52beE+woGUZivmROyED0vXJDTghchUHpQ+e17YO5KtpRFxsSUHa
0RKQJHWusvjgMbQrwYorrfAD+RHBEFFG+xof3NXR0R76+XwMQhTd3Rw4KNwXKe6PKtpFyH3ovKWw
oDxaVJXO6ingEqHPqYOIurAiuVRNEIEHPFk9+BZ457XdmCWA6g2amgyKQiJF+6OYhOaFLlSZZrOi
YzVAMmHd2AQAHquBLsKCH3H7Ir+9BCI/Y/jmiZusBBX2ginFBRdaGSaj2g09lAcbjvePyQM+k2Jn
9WvGPR3grQokoDZRufRaj0VMyEBOp+yZbODNj/ThL2pzNwEaaBCGDGwBqdEQlbmajYZN1VXTfhiY
lTXt8skn9ixXwHfASxvNiCcqDVuBIKclFsp9ihhFa98C78OMaNMoy88wjIszse9Xf9Y4lt/I4Fcf
C/ZsvFEuzdIQRzFa72tx/qQUcD1j1K6iNlP8YCNXMR6bvhE3ww5SeWBRNuWAIMa6LraCdprq7CXk
pGyZ7QcdLwzeC7ekl9gd0FjTdJRZo2/5gu/oe0CNnfDu8MHERN276CvhOzPWu/5h0RXMWXyvhvc1
EO01lxJR/g8Ql30j1D1SW/bReaMPrkqfPz2d4i+g1T7134uG/E6hlxOo5i+K9vfrtD22T/Pa2vYo
pMR+0PmdZxGTCMFKXjqPQo37ANUcTGUZPw6sg0jQVTqacf8uHoGO1f07QB6sYeR3W7Bpi1aYyZfV
bbXS5fF29G+7clZpCeSTM7Sy8R6o2uRGpz6ELf1ieLsdMoLML6u397+yLnt689F16KYyO0UZTdYi
UUIRIzv24TPYuqEe3QyzM0rdF3gcOOOmU2Ppo+ek5I0baoxfoTUVTflEdXKkJ73SnTaE3iVEmuTH
Rd8vEEfMHPrarlnICyWYxq24IcO/qAXq9SWs8bloH3idKz2oZUh0B/vFEQDOd1jVoFX87GKb+9rd
oFHL9ywbGlcA1mJxz+9gU6/yv59HpUrX+KHZAhc0AbLzckGtnTtkbk08ZYf29Ij2dSjie0MGVMQv
CvlB2BwzgbbOZkR2m6e0DuVtl8V1pnNhFoU0l03wFuEqgekIC/nxuBQcDGmQBM/RMWub6CfYpyAK
5y9H83vzPbswzUOUBRCBUaBmVAkkcZYo54dkgpGER/bjoFk4AQ4uksY/fZbiPcU61BGYp9fwQtJh
uPV9tk8q+BW5njhox1b23YGTPqGM4ZSnf4T/z4zvDPoHbJ65xcLGjBqor7/7P5cUSRZQo0EoVA/G
fl49QTn9EQ/Nifwvmb0s3xnFNL19gcD6erFUQN9z3ZIMB4ITBFI+0kBM6XkCCrH20FBeypSeJqUK
RClXOt+nAbD2DZZqt0DH+LXRCtG9YP37sR9SnTtYG1DUCx91u0NfUH7fNNlluS2GJP77IXfaGhbr
ICbJ7RY2rZok0bcp9ULO0lWi9Gs1avJ0gCdq/DzBbSSv2I9zWGqt3wTXYorwQRl/6kZ3ur2fWDCL
nUgiOBwtdxanWzZsy+EBjvJ/3bnIKnVV5UD9MqzyPrOI4FZcpSDZt0mfoWSIQYXUlROwrt/XzCHz
e7jWN19K3bXdG2WZNLvSoH9LFgfn+63i6bZhyD4ylXSkK9+sEVGLAweQ2sp8kOVxkyWGaQPZRG6o
bty0KqjLJq9b5WZx8r6j2B3hgO7L+EOv5w2TEDKvna/ZE4EJJYMz8SA/pGEN1ZnclQm5V7Uo4H8o
Wu/tJi4oUcuvF8S943MNN/LuLbt3k4m4NoPVXR/VoyV16xbUhKlC00jwMq4HsoErtDn/dbx8hzRm
cwKTfeHfWhms88Xxm57To3Pof2C4Dl0wqZSbmoE8Wo0e6XqxtwOMta8GcV3hIGhQkqWLtki308Z8
fpQuCw4xkEFPXL1uhaMiYt60vqQNFVEiEA8c+uJwKQmG0VBAVFxXiuVPYsxVGMhsU6lMDZIqDNkB
3JQUn8GCN80IUsvTDkv2AxhHijjV7Vq8yYYjwcEXDMzpm8Y8nsSKhgYPtDFL6uLlwWuGLtNCo+O9
7bxcf/dtVXHPSMs+7sHqPpnqtkwJi0ltOUKToxd9mmj7o0fvGWfePmyiarnfbqxGuuvgWolzlmA5
c7gBvG1T68XAP96ZS/MZtkuuLHOHuvVSsBk/LG+Q5I26ufcvwn6tpPuJkJE+7uthqFddADHbvuz0
CqlObrXCDBU7DfG5d4g9tHY0qYSTBySfkBXkrCVVEo/xt7LjCMO71NAWIs0yF97RDu7aonumGfaT
sNa95cGeVT4nHLwqp1U0PDiNyTsYb6XlsagOY3gEyA+9dSTZ+73FYfhOoz9HPE+vInHpsAGKJknR
wqIKuAbrGXhm8lzSDs3JWxW/tKHnfMnMNVw9dEkaz3OVJl5TEEho5glhAfynt8XXW0B7um4ZapTw
aFMreF9goQgkciLWomT5rs0lhrLBBTWS8ez2dPes+tGnwIijaydNr78zzPZGB35T1My/OBiC1uH8
1xDTmvbNWT4w0uK4Y1yn/A8dU6B7ETvHJP5Jxr1QW1lD2unzRvHkVanxy1xRY2clRvj9kHVqlFbZ
iJ7LnNBOtPrbfu+tzrFe7/ZU0Gw3qWrkm0LQNB8/3G2Uv5ePHThhi57aYhmA2ZXQ7492N8bV2p4M
dv60YBScNueG1MJKRLXQqtrS55w5/FvotybHkLJsUe+c8//ATOu0PlLhxYWNFB9tVJQ7mcyNsUWz
5dwzQgr1nWwFsA2CoODKZjyJNdkUuuGJr7A/cqc3No0v4Xh+XHGDBlnb3Lfn1KyLDz7P0DpLwjXD
2PG5/LA7G/Lt6g8Ewx365zLa7kpkmHTURzuTvgYqfRSMrR1fA2VLRsve6vsTUrZjpwuvCY9pqOBS
K0+33BiQqZl1oIGbqEJoppZ8X90xR+dTlsB1MXeDJEoxJc5fAzqtsJiMI4OqIU8jbVevU8grBbDb
2FMALkKwRrYNvOE01qoY3TfshR0AkJ2mWCE5kFcu5BF7lVOHZr1X7MfKC1V+/1SWspjcxMA9x2/H
9w2GTp7LH4lVPbKzCkpopPW5yhHASnoqt45KWVtG5WHWV92EfRYkgQmUq7OUnapZwt8yBr3gkVgT
dgeb7Zn5wC+K1b8Whr6zqdIzvQ3cNmuJvvxBr3OZ6sUZzeveijUkGQdAqsqQNLW/FhTFn1ir84rw
dq2G6zEAg2fpzN65pZhJHzmK2JmE1HcvGJjci+lPHjOy4SadVTibtdCKz6Lph8Se4/xmByG5Db4F
dKSD71DGJZ8ip0rebLbOF1RgaP+NiuMKSrtnTXZj4TJUyo4WdujuV9Xn0jyS8UvHOUUWKziRBPvB
B9cVo4IYnx+6Qzt8xNAuUwHn+ME9UEdsJPA+TbvkTLAPlsp/I57QKpgPBihLu/ItpC5r9K9RGnkd
reYlvZtJvaGxdM5dwO4r7r5xzFuPjZxvqErevGIAlHiqe9L4IzDP7jisBHGBYt9ut0oA00F4VrIN
ecv8ZJQaGiP3Zo7xjYYu4b3ujJ6qyERjme6eawRwYU4aSAHCIiZ9bQvgEuaXyFHemmAjUfHF1ii2
7z3f4LuCKvc84Li8S4vT5s8IwWIBBdlcL4Fpb48ZMGhUSGOCzPP1nnGIACcF9y6/+zNdFEpvPHCp
ZpqI3e9Q5em9Z3CE9v2P8uZ1qZdYx6LwTjn3lCNMFP/ZTfuJLqMRpsCFiEq+yknVPFoPIKbb5Kf/
t/B+U0X7RdDtehKsaoP3qBbTXVgfOap8iND4fSYRj3a9QzruFTOX0/HqTPIdjOz9BuGy2e7wG8Eo
ZvAh4hikbxDEdEJsN52KfoY4qRwwpbBKEpWDviw7VIDh7+Z8da7WyZ/a5aL0FOHEpjxSeeL6Tzkx
OBdeYqdqvsRnjMDZ8kU8bY9HUWdI3n+zvS/CoJhD/YTR99m0UKsvszdJBT1ioAQduEAlS1OIgrza
H2gKI6Ct6O65iUFfphQbDmqOlHHU5wEKErLhlK+mCqgx7i7PCMf3p7ZNEfVNnFRqmOZL0010Tpxb
D3rLRFvs0bzsQXQ+7SVaV5D1lPnO2RQj5F7OGAjRp6pPPKMYhlbbr311DhDJSWu+aNufTy/mqUI2
WSBmY04tMZuQ/PzS6PaI6hB9VpUvgzhvpojJQYZPC23xBK6nYwg6rEUcO/33Ig47MstHVc8RIaXf
1LPkh4KjxVYo09ZODu08bCTwzN9Ib15sR280sUPj99Lu4NlcErkatTNixMCdCyCFp5dmVVXpN4GN
AGZkB/BWfBXaxHqgKdm7KhMQW29lIEU5inacLgcqq8uGQPztKz5bqHLC9DvRwGBMrlQIk7uB7En6
OPANx5jvGEj/AtzDcyPBhu+NsihM5DpM97NCdbm7HjT4jI0tS3FAJlbpqwqYKyya/GpIRcaRfl5J
QOCEUdxjgi2qOZA3dGxuOmIYbjLOPc7EEbfx9HAt0Em/T1e7mecugp0UIBTI5qN4CD4pN9K0Aymf
0FNlq53eWmHFZJrvFN3j9bbOZedt7X9EmbAFrFhZ7RB2uil7xyVjMSHOsqp3LI0AOjJY9A9vQLGb
6ms6kaoSthtegirWSrKwc4Bjj4HuJe2xiKYwqC5GMPkkU0eDr+jtEivZaXzSONK/aqZBD2AR1S6v
9RIPTXDQ9utqIjRei8NjjKKbckZgDrIOgFTR9nvdmOxlCy3Ysdo4M5WDue1jmadr70Eo3BdbJiaN
gKM165NFH1wAJnuO7F/og3KtJVvg0rX/lPiRchaj5Mp6n4GvME649rSIbByiJFS1JD21LjhsAkH1
P8UOSyy0R1tdkfMM9veueDjt4bVBXyLxPLt5LytmE6lSfNVu/LryG7LzlAW06SvkuEkhnkt0CVww
U8ezpiSboicXc4ujtol3Ttue1ZwDyMqEoSCEDfetswRxsr/O1TKxZ7tRYPa/Zh9pmiqja2/r+urV
ER6gbAU7Bc4aoxscZgunymC6BWr6A2D/5mOuctzmoeGkmqjQtJVuw/c5SfWtCjsbZBqxiYxOM58M
DIL6rAWE030Zw9rsdlc5zbNLBMAoKI/YtIZslelnmvAij+DRePUjIVSs5qgz/a00DYdxHjsJtde9
U41a7Uf6y92XOS7B7UJI0+K/CGFYhCD+xxECeeq2KvdoNxwiKy05tX6eZ6EOw+V9lHEaFyJ1u0jC
Vwrr59McDWyn0K6yrjtv/hT7nAXc5qUPFEwCSPbstsT6bwphl+wUQaG4bLsacMq+a9+V9aLlCcgt
AArruU2vgG4CGbryH2lNaAU0l963/HuPUpCKR9a6wa7F+lonnXn+JzUsnBHpZj1tXp8JAm6fgxAo
ptUDhdw1vv1plB8V1UrHuS5OJImUKYEtQq3QncO/cmH0bTX/FK/gHYHBY7b97TiE3wNvdWUyKL9M
R+yxEbRaiQFkef1Af4i1HfleNpPS+GcAjrnn1LJ6HRgKTcsn3MbhJqOuCJlt64otLu9M3dbQ+T+J
32XoLjI6SsTFXEYKmS1T91RI6wjoihwkkBf+/2QYM7e2a/mXKn4HxTBE/pO3qXkYJRFdXVueYawB
0wbXJUlD6VqaA4LD1hWO24M+V7OewOiFpZ8/LoNqPk1nnZ+g/z15XEihMqHILdbt3EXLMcJwezXe
PcCHV3Qif7S4A0pZQRSOjPd6Tqc3v4xH8jQ90a306Pjdvytu5ynVDGkQ5kFg3X8xe9yZE3kfc8qv
PVb7UWrLLs246zjxBN8kfGPxSTxUVjMVuTm9OdaPdfvAxnQukyiLjD5mBrMjRbpZjzBxwUo9zhkI
WWx92Erp+FeNh6m4yUG6IJPF1DANfrsfI6YFq6Juh7TeiBrzICQuWEbA6FWMPqUvki74zyrWpyKu
Q7A4FslLPB9bWw28C6oXBcZlEat/4MqzoUKB1tO+ofC5ICwpGC9TPssFHvMxjPQ/H52e/TnblKx+
NOH8Gh1Ns9Sbt3S1L+0ouET+vkeg25gS8pgApba8YVTLi0WJqtPn1rjlfv3RT6nWfB2uPXZSo36A
L4fGrNWcNyLR9RpJ6DTUa1RjmRHCAMSggZHvnPHaKEYpRLYGG31J9pcXbikWqdlR537LfwE5FxTa
vO1nvWBPceIkaMr5USH09cs6iDb3TijL5b/jXqLFKmynvlneiNsxFSV2rIGsNWjhCCZnj+EX5fhn
Ox3coOZPAXv8IhkLpJdFXCaEz4spI0xwWoHmjwdcko2GeF0LrWg/oK6UNp7/ZW7noZGMO1M9yvN/
rR9k75MN8iPY0jm+zaxELcCY37yu52sUmFeBTX6rjuexR2F2TpWQ66E5TlcB+W7V9fsT6+mZOSZ3
8R/ILYynPwhu9OtAkHrg4l+bl7/rTIMicQcLXwmFJscHtsw8pwKpq/mqnd67/ycmJ6o75iw4tLLR
1E1I0zCpYFVBsn2Id7ib8T4fMhO9zuSbxdIolQUyWbmlkWITWqDMx24i58lOTteN+T6JA3KIJgNK
TrXu54XVE1Hr7QnvGGW1kDCmcFnu99fRpn62DajgasvJTxLcUbZ0A4sVxE0QGHA8mDYLHgabx9gf
bM78MEiERNH8sd3BNpiB4I5IDJALZJD4rGwM4o9/TdTzn97w+3whlL+ckq7Q1+0W4h1yyqFrKHdg
7H3esFX2DVPSQiqKXALqZliUOJK8xJ+OtAgaZEuG7fJwaKhzyWZZGCb75Vn5ejNprJoS6l5pZf5H
INDhmZzVnXxxESXvFECf4i1DC9/SM7p0UFA/abkRqc+SvM6oYuwZYgQOhfvSCIEI8d8GTngAltvI
f4VVapI9RRB0TrqiusKkEICTwFVR1RyjGvUZKJJXDiEQgaCJUDShjBWV/xgWBk9Mv+HckQke93Lm
YLiN+i5BhNgct7vASf+Z+3po2/5eY1Vq76x1pUAvJWVS1d03j8hPNlKDO/+ZnaY6WZ4gfCgdaNsd
y1huSQVwatvPopMKdv5r3QAMtQ61Tr+8gxHMf7JodtZyisDtIgUYpTnVka7+0S5Fg+n/BLtPDbFS
qgfdt7fW4lAaVyBqR002oLGICO+zWpyrr0e9T18zle4Ry2BdfUHd8aXe2UpYq1qALMij+YYqw4Sa
KEZvk6LjRmoC8QMKclKrmX5im7BUdlaz33b499XaPtUC+YWe24Vkw9rl4EXx4645lUV0S2L8ulZ/
bHOsLvEviaDuCF4o0iQLyry2c+mtBVVGoG5dtD02zF1BSbh4VMGVOCtIIbghwe5b0rGBbuAzk9HQ
D2MDD6HYjAEsgDoD4IaqujLEXPkL74hiH348+xZN2OzLDkVJQMn9zRLjph3Z9CepSQpYf43zw93s
aMH5S8Rgm6d5pNlX8HSFfNbKhStQvmeRWz+NpTjwnHNFQYpys25fzWWmdi4hKVijtSRH+JJKW43M
57cTJkhD4RAB86cHvUVd+jpx2vSuUcFnKpK6laNWyiK6vp8CGZzxo3qJSOf7xmODcVSGOwP0MKW0
c7Mg8AyDakE8qcVDsZFS1o2DJEb/dyx9r3Ss+1Naw6/ngvgsJfilBXr/7BJWZdN7ciMCtKTgx4Fl
bzhLI/lWmLLFHBTz6U5/e1wrWGc/+lgj1PXEQ2w1fR1b06tPyMKs+t2RIOouHKCxIU3B8v+myDAX
6bHVwLKm58rOro3zbFqRG9L/FnaDTCbAIyHZJEEo/nWXRDYSRV/zbjR1j0Jl1oJ7J/S3aDFwjLKL
7rEaKMCt1bCVqlYleyAZvEcBjukKZTKdIQoC/akwJFMZj7Ev+A+7Hzyv3s1VRKNeMaW5hVJIDqBE
aw6KlhZpGYkBQH5y63HICVpY8KHA8YBCFW9bDSNOus1HQljdy72EnAnTY7yl4Lwsq31wnLtpLkFq
Bv6xuaF8Mvve1f4CR4N/xanJ0haDAXX2WTdSFCAEvyqPMbRpJEuj1sIsdbj6X3qUfegAKwDQognG
d3Y5HlhPlbrqDXcVfaYfDXTLjhMJo/Q0KEany+2bPBo7IDCcISwONrzPtEsZlBL4zRKmmwqfU4bW
miwgBhF92cx/WhEDGk9wL5pI22LU59RT6VIfFqUOliHJW8o8fCMpWbczi7D7jTEI4LF2yUUjSTqS
Mw4XoL7744lnoaeHLCX/EJiJ+p2tA4jiv4kbN5QjL8ujwAHmroDl+Fb3p//kcB8iOZaXIGQAhEwb
Oy1xhbxrT8ZKLwI/HH5AbsXARnaF5RzxR55pSBVN9LZqpKkZvHFugy2VdC2UJJk/pYtWehi+bnoE
a5brvAK7MulkYC4CirY7JjTgHVV5/etOjya+nJmNkiv/PRgxdXEzr5vTCdUJuxSJcf1SB4tI+unn
x1aFUh9sy9BUvxXBgCOp/OYjh0pnpbDPaqsaUazcIRsYdv56mwUAFx64BMpCF5sqDqwxKq4oki1T
rVVSD+G1WA1R/1ILF8DYye7Lfz9N/0JWrov8U4qOrEKJWrtWekwWzTDtJGNdszW8OlZ5QnLDw0G6
UgGpOov5NBm0OQkG8UQlIUPtkO4gvD6urEfY6fz7d3wMkxiGqPNqMAaCNxOUrqaKCrvN6+plAtaZ
+bvZcd2/C+pkXFHYXRZ3MZ9K56klbd+yNQctZPGd/KkoqsFclQZQLRsarT1drO/iktw8voaQDKyq
1KKqPQLzahGOrRV0+31f6IclzLeh7yi2Nu+ipMNV1NDQvsOrSdKNoCY0ZVmxi53qyRAULjNDO+K6
xUj3PNtTbANWw6qx/rhdsRXudPtGFVI7rjcUpuJKjNgYzQI5r5eHG2tR7DLVRhzc5ju5S61pXv5H
0Z0uSDGmlbKYoKp8WXkv8HgRxnKvSY7oXL5zu0r5aaGSsLFCGmgeCOaD8VkqS5aybCBn42Y7rNoN
vM0yWj9sVOSaHgRcEwSeedn4hDNZ3frzcZPRPsDp06nJdQXVFwmSYEhDQTm+3LX7x41Bj1E0tbsa
uIHxNIjyZ6vx2CfGcawvqceXCvGwVFOHG0Ftgw5zSbeS9B7fwKcuSzsbd6xkAWx7F6gzcK+6aolR
iEpMk+ygWQR5Z8rTjOGHyQ32dipn4YT+bI2tJhadrfYuWT59kz60dBo4/mRsDwHks8OKBEbiJDJR
0Q9OXR2GZ7FS2vwZOSubDDMkTAFJiW7YQrWV5UvVR0lw443rddqGgDFRaeyjt8CaOSIjAp7NkVe+
3YnaoGKqfo7MNrj81I3/ynNc+xh12J90AR4oj57KZv2mCRIzLBBXIWfQEXKg9EbzIR9YT3oMsefu
0Vr6i9G7xo+PAqnj24TdE8Btb+dz/PR0KGFx2QC3Zx8VEdkrZIbp8Ll4JseXMLrDrv/WT7EHpcUG
cs3BPblWstcl/w9OcPrwlUqzuZvAYFzPlZ65JkOD/nVXAqnrPIItwuTVP46IuXEme70WeT+U/7WM
M4ylisblGkOK+R0N5y8MkMQNwy6CfJKJtdoJFxRT8rPRx8WHf0Sge6VsCLa4zL7fIfbTGajOufN1
pejSwd9RH6thhdx6jkMfxCfHxEnrohP9wex5DpGyeWPWbm6y8XwDzVk1D6TqGvgAXpZiCIxgvnGm
R0ClGe0jjVCPgPTcpn/7cjw7Sd0lBy3Dp2VEHrHfZZHFdm9Jnej/PUSZyrusMoTrNgPJnUB0uZHN
jG+nh7uk0hr8RbVi00nmlce0iNtUXAHDch46TLIha0j4llbA3ocVPRLG29zW61bGthiVUL536rPL
4gHkH2rqQd/+phSF289Pize9C4Lw6Iv606sx678/SOBdan5kbTs1cLhOHpG4TpuqEDYf5l5n5AUQ
pKSdYkDN1Uc4gtvT8WOPlLa1KxxksZSgdfDi1+5td+pw7iy24I4X0rRrl44VAT9sp+xhLhkdIupY
5Hei/RLDWyY6BLrfJgfSn30W7dNP2mJpJ4RiOzszjwB0K7uylTrcuXCFr1wIZ19wrCc0nYkHZIEr
kVLxQLl3JEgFOybhAn+chhyNjpS8d6IoXlePemICqUL61uNbQdPKqtMu/G4tH3/vTzwmNea55dLY
BG1NiLKukFNoEfKfGqLJV4XNV+nEyKwiIrpPlXJlXtgrhYOJ0CCOw1LB/39gqnjKQ+hvmOfe/oJ3
9nbH/ttSlGFXBFx8HOmUth7j9HYpRmkygD7p8G7GaEp+mF60YejEojYmBFN7X40CFtr3O7I8lDrb
L2eK6DAvfhFCpRdEVqoKTP2f3qGiOSjXGjmkidCMA5j17u0KL4rtFKZ5gru2fYUitgMF5D3ajuCw
9V7R8A9Igti92X9ZjZlEQUuHOL8UtnKTX5Lrt5J+H4vdi8mHj695NBbYkaNn/mVCCuGndZOYgKa4
SwrwazV+whdV9xo1syJ4CPEzVWZ5145SaSBXdkdgIzeNYTqxvLpbcNulwA+e2vfYMTZ+qO1NoIZh
aRxi9lEn7i5xGDcjGVKO5V6XmsKuA6ZfnoYuWl+BVqWYjFh2Bgdbg2yeJkYPsQogcyIEApUW/Ypl
csHKvqoDRf8DR+3FOFmKOs1bqG4xJ4TGCpeMkQhxE1efa7E6c0XXgfY05MtlwfCFsu9hNKnoLdmD
u9ydKFUpTKl9+Qc6DlFNJCjrDFyt6ua7JT1dgcEndZmQHCHR5nZZ8gYHnpCalOzU8m4eebfxQNG8
H4QOS0Zj2Pj4t5GvfrUnrpu1NVWCOu1hPNEMfScWqlcxdx53YlLWo32UC5RSHiEiW/uMN+VHtS3V
tozR0HSFGxw325DKV49VMDdxLtJBQWTkx2XtuYFXOdIJYUJAcXSTHQ1eM275u2hwY8LR195qjjO0
UE1pofivsH7RmO+yD4UZTlvsfS06kJ8J5ROXi86BP3e85D1NtJUs4pR/xHTCmcjev2Wd2TJs3gXw
wgDFYFKWd8Y1AaCw7g32VeCi4YIVRzWcSmTw2FH8MdKlC/KszeaBWEPzo8KyBazSQM34Gy0Nrf9w
ZLd25ZoGTJ+vsxNAVOxSgP55Pgl8KIY4T9uf8bv/e7FZTU/PgJcpHX5ZF8E+7QeXgSUyeNpt2nK6
EMC2il1kSdG8P4xQpn934ZYuWwmczczyhkPKgd0kUgqOx7VftLG11QeFoRRXaZ5fj0eeYvBvjIOS
iNvsCcuV22in3xdKk2qsJL4ONIOiBSAuoXvrlavvL5U4VByKqUiUnQvcOp4FoL9myN2T4sDqw1Vl
ndjhRpsO1U/BQTeK/ca9CzmNGrKYEp1GpACNnr6Uae+ecevMaCWPJUYc05SYNCx87rkq+Bxfru3S
QYehEDfINWnPq5iQowYoQv+7hi/eK8dhf7c7tZ4NQFMtCFRfbZ19GUDXOiW9qfhA4FcS5Pf1HoFV
3O4nOJjauCACrdObyso3NPOvXb610zAnRyxIaRGe1MUq3gonKmj+GX0XCXJILg9t1Y3ugowaeb2Q
riL82ZQSjEtS5VPhRL24hQX6yfxt+EOtPoWcOeMpeiZNDMoEM+iNkTYl/Fr7uIidB1S5+e+ppoYh
MWbWYagMJPLx/yuuQiLePEqhkx8uBtGDVfeFRyknEXNlBRdqalrLvhDFdkEo7/A0tPHjSFq8l4AM
crqXe7UA+gmzdfE6Z2Ecl0Aw9wLuqvwhVN8TFLcC+cXcBIYPRtslmXQA+tdylFHrRTOwnDWWH8k4
lgk1kRazFXe7ztZuhfHmL+8Htacj6pKuzSTndj+xKnOJW8Ay77tPKvI8jTMK+cD6daWMqUPxjfEm
1L2yfs2zObmB/uw6wI74yvfDRCLSTwUe9atA/ZOhJFywWXok6p2h/poZEC+t7SodGH2J+Z3aRaMj
+rtTcivPdgNMZOH5lSdAd98wLzfe/BGhlyn8GDxV1tHlf00K2xENcVITpIKT97iTvL9mKUAQbw1O
YHKQZwtxh3qBZvY2XkdbnDtMdB8PPUja3zpa+k38NM3G4I65pavdU5YcGBnsaAvhI7djl9dXXwam
Z8AOXiV0KALsdYfgE32KUa8W3/7aWulxfwnfstXXhRtupeWkJrdMD03nWGXyHSWU2hfJfkSnIvO1
I+JC15Geob/0iGToPUoGWKkkrfzhUbBb6bvNzzLpJgHxvb9YlDTsCP5ZOVr/BIyqT9zweU1xNLKI
0piU6oFi+6X7fsjEE/Lo1mOdXcidteSv1ecB3HMeSZZX+x55zi/jAxhIz5MnNjtDCSgucBpiUTE3
SrFBaT0Rvk5TRQ4jMxwM9gbq6JDDdTXWYlJDmFMV4b//zwmJod7SalRCb6QlKgb2IZlGijOtGY5N
3g1wbJPdO1ArhlI7XEDgF8Obi1BiUPaSzdGOenzioh2bJ2NQWuSGVcgZ9f6wCVr9aJ+qhLL7bfD8
+rd1CpOPut0Esv4leyLU5axph1jxdN3rujzkkFel7RHBX/ujodng6G6XLkeYqw1L5w4wCw44sQEN
H0IBCSUUNHygxV8pIHr0nsSI3HSY+n5FJwKiTw9GpoKiTjFhFi/N9o71dEpQ7kSgCumIt3ObCLeI
1s4B/UMviqekk66ox3BNIWcJSW0NFSmKoOpZdIOS7D++QVArcDIQBYadyXAw1Rhphv/J1XsHHnsy
U0hF/AmOH6yiCliGji6AhGDGKxeB6uuU1d+mh6b4DBgO7pPR8VHPSuJw1dZcPbIdsp7zzNQmy2Gu
ECpkqXsX4S3QaR44G/IzIt40teqDPm2OGDQIF8ICThtDxeR0A0jUvrgYGEIyW4AH1DxXVleuXswI
7gzxm+geuhP80vjN0JQNXipix8rsg+lwFPXuYMhMp434XkweZA5Lfv7UH5JuQXIjsEY6mf7jeIeA
Irn/hkdfGMUQbcPAW6GL/L1IN0WOUp+36dh/o/bjKyLOZXvojtgQIgt8WiJKw6ex1J1pkXdWsD2m
qnk7EOnrZo93RgIyIG9D2wv0CBX13r98OEgjU/mAQ8pRg33ACVyCuE8I6MVfy/JG4hXvAytewAKm
BDhresilYJ6Jm5lhxUgmUNm2At7i2T7LwWDdto5rWPsu6o28NdKAVDa8CwjgbdHnTF46JdiLk1Ah
6k11s6s6ZKnL78yzR7YSMkiSXA4s+nyKm6uPS1Zh5d4H1vGSj4fclHHe28H9r3dC79VNqBzM5i1p
XjHt/3wzeq6ZzmmaAs9pcv8Sper20i0s9sQHrIcSo+EuMzYJS2RbpSUCAV9N2l5fc8EwXL51EU8J
CW4yoQdOueQ1LxUcFIYbeDbkV5EBn4AmbSeEKs7rVof7b0/MLiplwLRmGeV2FfqWW7HpKW/iTWCf
VDwwv/TpfXZbuKVdy0iJGzu3Vm0v9dXw7UcU+clI99xKoVLL6XqfSz3yNaOo7k1h9ATK/rLuE4VI
X7G/4oImbPIhcD4cJEzo+a+oqA9i/c5mCVGhJ1r18bhex5s0tWJh6HRotRRE8qtGw1TabA3OoLQX
cHcJgWjdLEk6IbPuf12JprOiEU6gQ2AiampsszxfmK1S8SHrK4tO6qPD7eIy8xNSMUrXmtWyaWZw
4U4pAsEJuF/9zFNhD2J+CA7cK+45FYlldcnhv8LchYkL2bV3o8J4t2WjsKQNVzL8Tdzn83XSG4YI
wHcXlQblHvbZJFwm1hSK6LbWOyE6UEzZHOO401+FKaaOO+Ml38yodUnO3ZGKrKfbFuHokL6lK6mr
sDNqhfBh3tbTvH9/CfkWo75xJ+mERWMDS5itzgOvqhH3gNjoJ8NW+Czohr54d2G6TK5zTW56Ndse
TLGcNZthm2VGt4USG35jjag2RfRZ0BLI6o5ghz3y54FL3RwsD2OMz/9nf4k3xfyoTuF3IQ10Wkk5
S9daJJQSWSSlUoDlu2UMlAqqTD/caRkmc4g6H2gC6g0G6WfVFjunguhU5Mnd76rzH1Bjs6bcE0gD
YKhd1jDBvnrRG4wONb5ZefiZo8rFTtm85vZyiH5uOxvGS6xpS6qzbDoNY5VA0bVn07Lw3Z3YQJe0
m/W+mXcE8aafgktSVK+F4yf8DlBZR7up88a7OTNom88fgpwuqxjWkKbC62H+RDINch2eb/YRWMuo
kIFoPE0vCkGTZP6a2egD5eRDkaw88GrzRb4Njnd2pGPN68Uv8cgEb1v+9YKMUzzeXmJyigoZsTsN
KDcfezQ7zepVyPLF6rdRfmq16VO/Aueu7E1FgGfBlkDsClwQ03c4GPVcgL2af4eW4c8YCWYOSK9S
UU262U0YTWRUf7ne55dBqym1HkhmziIj7twqcsJRm/vjlQyX6oIRwDkHY+1AVpL80g8qExNX2/gc
LPtSkE2XEwECHsqGRSrOeP+WR862eQD0iSbKP0Lm0eC5cMj5Appw7pG5RX5wV2Fo0vvuteDTpkmk
aYZx2nXpD3bi2jD7ijjMa+rjxqeL/+AvujM7+RsCMHPT37Acc+G1L+ICJ5LEYbk+7M3fiDGISqSQ
K/nzuan798vIJgaPoygE1tDigssvKLeujA6ZXHeQNvgamK7r73/G5gzRkA6JjJ2nre1fVd1n9XJ1
YAa/LLcWfW6vnGVCV9QzwgTFzck2hW2RtrkN6zxV5GViItMsG13tPfI5thKbyYEp+rxjEjHA/o2T
bM+P2nZWrVrDuOrTBF2jmmV4cumrekcWv1wJ6ekRpszJWSJIU0bLPzXszUSFQfycnw7iIfa6lcXc
mVSQ48IA9wJgZphdx7hOsES/L1lR1dqsEgH1J4MlEohSlNCCwwlifObBO4+mnDllNP19JOGN6Hwh
jCyzZeM8CpfaSsMGUYNUZ3citvat62krN5K0GdYT09xdZd9O+788mCfz3o7YK81xjybS9Xun6cqV
nEJOBsdX24EcxN/Dp+T5IWvbHxbmXuM1QllKUTCkfskooQJY/w1/+p9FmyRtlL9X6nsQIuIytfmp
XGE7ccJ4A540ha+Jb6rTRto2g06LDn/N/MshhwPBxBWelB74ynWEZbr2qdgwbpu6hfWKye9f2FMN
RyFqrkffTEJr2PLdypXgEJ8wkUdGAmETueBpJNScmgajv/c+p7FjWcVt2JyQDn4X/raTzaDygDX5
B9UYClf2x3cTmyQKP6yF79xPGuTLSgKh8cB7okOej+Zler43zmEEprP1JN7qPktiy2x07W63gzOC
bTxhLMcUX9pNVUGW+tWhrNdmMguNPjZzSHJgA7/hnouHuuzI3falOqzD5GEq/jNRfba7fWSydTEO
SbnU8XepgGjWJmRezdogIbOjj0ZN8Wg9Jsu9EJsTlZL11dRUm1G/EWZGGC/vYquxrTvoo2zF/WOS
wnq/F/OBLypUtKKqnFDDsqIL7bi6vaa/yB/PmmO3Rl/2d4eMDZX2j37+VlANoyVL9bujfB7+Dh0g
mM7j64vb2UQy2oIz+emXk6icIIl1ueQ6RzrMKd7cforXhHqFDddcUCbe16nedm9kLeW+DR3I3FlS
WPwBUMGQLQ4Xj2nUMC62ArGlbm2+E5urYrXDcF3Ig00zFWW1Ubcg/H3cqoEIdYO/FKSymwvnB4QZ
kAs4oV7N3WtzbMhgML6CdophpBnINHBT9/Q1r+mtXKbMRLgIc9m717hg3oWqAZlvkgjnZ2Oh6QVQ
YQkY3DtLIR+6VMi6JZwQ99RwEattlp/2kFzRtPr7wnUTIHtLbdG2SPcIzSRqC8G68nTAp4J8QBSf
9lYfGWUQwnjFdt1OV5vU5YKuG0x79zhn54pRIrmSZice+Dg2+9Y4llipJ/4XCWpi6AB8UdW/coYE
1zsfSMLUQDVhfWrxX1RFn/wGrDfxGBSM0sUN++gccZnUZMKpfuzV0nqlyD30y+552B0YQt62UjFV
TBWJhDRw5KAILVGuY8710X1mrcSmJvr3CCS/4cEn5f0Ou+NnLqst/0frpUJT3jV23LI967yaN5B+
FmgcrhXLcnGkjncwV7TacYjTxvp0A1kGUNRdaZiFTXUceUudYz4hVxPDYmppop1AnHXoU45etaND
pG9VkSlrYRNGsO2j4zWoE9yq/dYaw/mYr8e8u5sVGVZounr/aHzD7CLGvSoXn9a8IvB7G7FEyymR
1DCv2fj81LdODmQLiJTopm0vSSB0g0rqXqRAX+uk+sEgOere4Bmw02F8Y22Z4JXjKDZHBT+X4keu
HNnSsIBegIB/FRIQc1cBl8/TIyDRNs/CagTXq3WZ8gGNzQivEq3uHBTgjHcDfrA8YVxZ40o9HQSF
UzaOPof0aKJ2r+lkDg7XxG56v4mgvo4pfliOpb8DETqT+3lPL4JLP6uqt77BMp3EDwZzWi3sGyNE
Zjn3ehFiELJbClj7lniIwY5Xd4mkjm3r13I/8BSXtqJ2M+8HRmdI09pd5W8OqXWJPMAYvTizug0F
Bopi7505Bdztf6BM8+UYTc5WqHHXxkBRBv6BTVJUggxUQacezuRhnrMbW0YCi7gTbzTZDE1sb+17
yXTWRtbOUETj4wO7htWLuG2xhhSu8rnITspbq1DE94+3aEh4K4RJ5XCPyPRsZFacLbDoBQgsbIA5
4b1n0n2HfS85gIKdgKYFxyMdk6x6kWcgJ6o8plOMsxBYw500oTF4kpwz1LIIICNGTcr1gi30zNGU
56RPbUC7ydR/islzqbAO3XTp9T8Nso4XCB131DcZFvJpciSaAcBxSrtTdkNrC1LLXWEEv9keD5+D
ynFwCkSRey2DKZkuLvV2UczC7kR2TfqUfae9qw6YGzkjgPiBGidWShsAC3EpjOlMlqW3QRH0qNLN
doA1GSZCFA9CAjCxNQah7VY1apjq34X+2KhsKMrMpEHZ/wfUNfALnIg9RA7j7SD+hWSH4rlQ8x97
hyE5hhs9LZTAOu0s/uktLZ2Q0BbirDhUFGcUHn7d5fq4H8tZx6AZgNq+1aZkgGS/jeGc+84EEa6P
2M4bJmQAK4IcgYYfZ7xX3exQPlRRUFHoHO0EfjeO4Uq6bMlMA+KnbrtORjsg8Ynn2PttHHDtX1Uy
lbLGTZD0fNs8MIFWmTOgZJoeB9jUpInfxlbf4JjwyWiZ2J3/hreuclNG1vFllPNWxhDNqh+AhTVc
gPTtkhxINb2tZWLeuufKrwC/SicOGMV6EH/Wh8u28XZvR1QAgJWVGvdYDrMl4TdL6z/Xxy2BIZFS
ktTaLVfBbXn9CW4CO3Ol1gy9aY0Sgie4idNBOIsKqiYvWfhqwszhlLh6lAQdJV4yXRPO84apOUub
9v9J+Bi3oSYWvOIGqWfDa8XYoVl4L99hvyYUlcKYd2Wc5oHx8ZdbLz/kzBcFuqIDeZWdPYnaEqVQ
LQNXxKcih06cr63mzDk7icWtLySollPtxEgPQuLVNh+upH3IqnvHIsM4ZHn4J1h1M4siebt1/dcp
Ul25fKD5ZNmOAaoeVtPy7tRWwbb1a+7d7G9SNUkFobI2etARmom/uxyPHHaoOAo8bPDUbLLZprq4
ea3Y9Ep4oGEkC2OfQnc5AtLsFoK1n3EKIgAxNZYU5i5QV6X+aEGDp0OXtZQkdPd/sjrhBd853+iy
wKjqcQXKbB7My4vQIM121znAvCZBB0FSH5hTFOprTjyJsn3384rlNEkOcOGpjn32+gy+ZrgQpujl
1Xx+GuYctzbB02suMY7BMZiYquSoB9eznzLonrUm2lVkWtukmSywDPChTdV9rctQ1DQhKaJdRwI1
G/qwrQMtv2Khh9IpP/j6Ym75m301wSwmVkk+aZLW59AFt07baMKuArLsodf3j6DxjSA805Go/eT5
wDD1hwAuxJC7QK/NprtpbdwYsf2VOUXph5K92X6P3ZP/0EbOyWK8uzqsqljTrXzlfY8o7pOzoeIe
O7YY3t+Cbqfr1DC72utxcxlBQ7qQAiSruklMQdKoxjQMhN77zn4KsxOheAz3k2fZGSRJjHzdLGbM
s5i7DiNGM9En6Dji+h9ZbLdSVx5VVkimsKp3sqoGNqm53S2tNWB8u/nOlWhZMLAl5vw8Lrw1AhF2
FEWAwrqAywGdWooIP2RTUDe9CoVkbRyaCpEBUylwhJYOKW0wnAQ9q0aPPLwQmBejqHOkLSeK3yoK
rrsOLWxj/eiZarnSaAerLLd+bELAGbdLc/1MM5mFHbty38mqDFPqDKxTP0t3qiuMWwlKk19soe7z
NgtNh7VuB+aMsb4wHVj53rl+N/S2/X//+23ucFS6Nrv3YfL/R+r4QCmo2XZbRYc9wCM58K58quE5
bdlyjR0gSOmMnODtRl9b6ZdhYAe5xZ8ZFVB6RQQpG+ZC+3WEogy9IoFg5fVRg4kfRuqrGHomw1yW
PWKGj+sPtj0Ray/URQBxXYjZ03oVsE8sALZd9/zvX1itc1gEDscp4J7Cnh1jKocaXX2sm8d0wd5a
e+vtTRVTWfsHb+NchsnibwO0mpTYiy4f6pjRhoI34yNgJmukMopAu3EX/rvgndO0i6cXvRlPNzOo
aoPjTDh//fukH88J9nDLeYh5CKZUg8gJwcX6c02SFbyNTMM1f6n5zhRTUCmPi0otrKz7ar9YyrsQ
sOP3f6c6FLjLiAMC4glsbVPfogcRU0YnimGnra9Rn6yRxmNZiKYqcslaQXBxE2ykG2JROH9DuzQq
XTrS1mKfgL0w73N1aNndSuOucvtctEDte0JGyKiDqpxd/FAOhZk1WNVn8ahc3DjLJT6VB3kb9cuc
WWgs+nm+3+TmbCcAPWZvmL3ug+HakB+PiozdNc6WJ0XTqJtBXoYaTStF9xZ4BL1VFMY5LKbX5u18
VNVKvoQ3jcC073ELp/olcfN21ZssYKrqrAHLnQ7OufEznX53s0BPu5kXUrvnC2qLNfRQWFUJ+o9e
xDTITihc1OGlcOJmvLHVRpALtjzz/cremFQxxrOK47mu49dZgXQ8UAVmZysr5swtkunne2bF1p4V
zcFUXec9RdsTMo/Tele+gxxuaidRjXDRV7dU+OKu+jIA5TvCm8SDZUuvbm5YDmergl/DcOE0EdCK
/OqUonsxLq6/6CSwnhz7whC61Q7elKiSHWg2MXlJydZL5Klpz0KRiH68XK22l9BTpmhAjpe/3nKl
cbCDDLyfMuMPOGJ1ZJPA9dxCSFc+SMw7rzYFHTESgo+UNOmiop+7Slr11bpVqC0hjlLvCrQyV/Gk
O07icY95byJr4gYgH9wN5lSo8APl7qC8EtAXE09JiQAnbyBPBjzDRSpHi7a5eV4bpMlWIWVvkiaS
EnqGgVJSdU6/r9g5XagVxOLgcXL0mnvGg9K9yA9O5IyVmhMEt4BV3idH57fqjBWbrDS+SpQWH7aJ
T+fqqHu43IQKZ/0HLLFpb9BthnqHox9vK/JQEfyV3rnixoZRVpUZSy++5cwtfVaIwMjZsEA0zowc
c+fwjQhR0RYRgH0s7PBazSm+fcJG+QHj9J92svyQ/7roCKNp7H9YA2llqPWTYYOvMQybuze63j+0
f922UMlZcdXTSFNYoFu1CU15u8Wc/0cRx+u1J/Wu2amInFW1qoCABgzSUnpQ4Tjd84Z/jQCpqyUv
0Nm04LpxXluRc4N9/URrem0l3+oQsh+XmdtGUMc+GdJyswSRku6/fXvMc40UmHIaSOuREBaleAD6
dZd/0uWRPBOs1LUuDRfzsIa3NeMJOfke23EsgchEp+BfwHAjbTYd8uj6OGOHkoAM6WaNcJu3VrQr
nd3FjLeh0k0SUIHk0OXjejBW8oHUHmyOnysE1vAj+49CuMlfJJ/8mykdmuLnsrwC0C6Ej2zKot5K
jBPEgDcj/DtMbsA9Flhhml4fLTtTB9vzqDLjScnmIaZDJ+SwrVJgqFte3c9DMSP/EclfXrMyUbHY
b4kXN6HGiiDpPDVGQfWEKqhWlQfqYD06bSORCflw/e123fjPoVWxes5lh0E0lMmLIfBEoge7mcFT
tOFum91KZc9Y8w4Jfrued3hTIoCBf3c+Z5P1yNVg9uNenAHhdofGml3lNIOzCt49cy5q58j4Otqi
JhyvFWjTry5B0EUdkNVz2JMLZJeSTjv115EDjpcNqgAeIJAy9SKKMZr5fhnV1wvbJuMZ0rffu6W8
kzzhiKza/QRsHYaXxhQ2D7IGQ6LCec+ibpRvbVzpwWKrNKSwGXpF5P4xmitAKT5sy02hlueP65CM
8ENJhNkIKUMAnCS91ZiO4bnnqCEcNOkz9nTJ0qkKvIQqFqiFQCkiD36I0jF44VLar3YyfaX6YSXD
9HQL7+eRAngpNPkMPOMIFctuEprmD3rfV4XmrYtPdqcudYQDurDq27WHk3PhEJg/UK+psyYVciX9
uSSnzHPypenwTWyRfNlb98Rl4Vw6gWnUKqwxoqy8l+73pf+0Zw3DskLl0yybu0me6T/WGq44EXkH
mCg/JzQ6MAkYqx9gV+w1wtWcF+Tj48RBVcXw7Qa3UjtR9Mc2li1v2jxgApPz1dnGj6cWsAFmqGFc
zjbR1CCfr7NxlJaJ1GdsRdKTukLS5sEE4jMMKWuSTekFUB4z+Akn8rQrRs6ChdQptoD40MemkNTB
py5VDYRWI/2z4E+1aCNy2rY1JMIssE6FJMNYfbPIez+dt9/Kt573EwqETsQm6NwPJaWCZK+aIgpc
DR6pj/WzHI+F67oBSdJH2YIZ8dcz/BuYiAtVyZQGDLLqyjDlJQTlpWzEXmcAVOzrqVh/1rGBvqxb
TOXmNCgLMYthj1/3ujow/qbEu1YWbecDqO+ZUFGOWZfDhIVnWokU9Vjy/+cpoacN1yGiEaRjocEk
7Q5fEHMcKbjoBkjYWUWxenT9y2bcLtw/YRJCuSSzTceGqvVPqfOHqtrrEAwMhY6EJx02kx6CLmEA
tIxWvqSfl+fVGemt+PiVGBfSBb/4Ev5uA5XNmFDf8kSSmbEgrnxUMuxInP3qZvUVSk+zn4w2D1Mo
r4WUW1JYFNgbCUQjl40oooOTkSiTE5dHCl9loutYAcvAq7ARPzuIMgoPSe5mIL2ewxmjd7AicoFY
TSsCYoYFVnSNKdiwXaw/52C/ttUOEE0ImhFd9DfRpvZgthJeA26zATVq267R7o20UoqwVqws5S5y
BuaSk+upVY1qMIf49ZT8pd5IKN6KJ00YNcmsXeYWg3HJJIhUyZ5O9L+JAQTlyBPgY/qRZEmSD8wo
FtDfu6WBaiqFo8veOwTmk9ozwZDKbiD30yiJmgxVdFHy9ELokKvjhlndxOIqKDtwUfTMvVTsMV5x
pje0nKndgh3Wm3rYGg8GOboUcpM0dZLSpmm6oJqW1swsACrJqqENDd79vzzeT/ODyZwc88ZDDNTv
v2xwV+2hfdVI5oxn8JP9vZ5bg+yjco8aGzc8rBl12u2EdCAmVTYQgQKx/+iExEy1kFq8ZD/DiKRz
VkmKSPWEUg1C4+gf070fZgfNdZ9V+WzyTpYTgLBKRVA4c2a9jho+MWVzBXwb5XNX6Md1gy6D0kT/
GxP4FTOf+iRMjlciUjUdzfp1BYJ+VAJLvkiMOUp9en5XyC3sC1mD5fVN5eEMvZCENzpDNW4eO//m
oNUAugShCrTpspgU5zu8r/KBQLmlk8R2f1wRUSL46ZFOzUqmdca0vMRK1JPd8qO1ldUx1N/9BFTa
8Xkx3w5JshXGGRHGk3qucKY9eQn2R/izg9Z41Nr4G7WGSkSF7HG92iRZf9mBuv7Z/c2hJ3DUv3kd
8dFiTJbYACKjcZZslaZp2xrptOvdeq7+NCxRczn7gG1+8gjXMKsn9Pb10WPugtlNlEx26XsqJCWq
Yeh3r3ep8hxI5573xp5mCfBjeMK0Ge3tB1B1nZtw8eRxI5krc+qfm5F8ZsjkdPGmASLChn5dgQY3
ohqZIWX/P/AHlBQyXdMU7ar2jV4CXTOmmJ15wk5TJgQ2ygnP9FPeX4fUxtlnksiiUCmpDs+nn4N1
MLsnH8y2QI2eoZM3wE7rimlNbQ4aHSmQOtN2s9yKr5dlmxSOJ4M3E9Mkn6TkiPGX1WHeHHuSCIuu
EHG8ChphqVYluKBvcaIbPcUowdAWLJJmLqxHNLEmb19jR0Ddvaz1dhSACOB0AeGRh1mfx9vagdrd
b4NKwDMlix62rAZitYcs2auQLZaRPka365txs2cHmkwAaUORjw3aKUGol3iccmbzE52T7nZEbjri
Tb/Pfe0TtvHR8bV4LF9J3mcdrRcDykkpuzDop/0hrzF5QH6sWKmv2Sr+27Fq1YY4BM3OOIPuVsfo
sTTJwg2m4BrESS8Pu8hyH8DcjZ4QT3koY9yJuPkIl8NNfsO3J68ykrt/cl/DqkvnSrOBNCorSHaN
c38vLsyjhxxgzn3lizhykBOOsjTBgMRp1bFZek6pqyIbrwkZnxf7Lu7CtMHefywSQodmzaWublem
F/1OQYKprHY/9HZJNpNf4v03Ou1QP9jvnOPP/oBosvbPtUptbsM1+dcuRc6ssmtu60ObmBZA3y4y
EAQnUnSLpaaC4Dc1/awFxVJZm3x4AzYCYez4+GgUQ7C6PStWDFlQuk8+Cs1lG2SwZYkj1H60CBN7
z4DF/p08XusgYM1fhO3RcWnAZ3ngjrG6A3bdEOvG6RHRBonCBOkBXvFkHQarGGsNCY13kvE1vsfH
PlwtYXjPgV05MIYTlve54EC6wedJgac82YnOU4s2Opdv6G/94hn2l8oO6EwD8gysXHByPBrsN4If
WQ2Z8dMeCmqDcQf2QsAkBwBDdjTdpL4xTarNehNz/WXrIydaLRBya+ZT+eGydh0ByyOE0l1CDbqO
8MGBI4xORGSAfuuP1s8Z5++CkmW2LUEmY8LPYXlOjE7pZ+nyW6Yqh4thpLRxCu13a2KVdPbnk/Ej
wT+y9lK70aCvtxq/LLkRW268hTmmkITZd3aRWBdFtnDWZ3ULuNle13xpAadyYcOqB1g9fBLEsaUg
kB0HGQNycHMX3IIVccXrqgnY97CmYgWa0IgBFuRY4Zhb8MXECH4GhPx5z+/AkSHoGNMQex/zBF6e
eLvSkAURtr3ACbldEjiEgtwUM89PpMcZ8zTxfdpwawPccx2RUgvvqa0R5cz+KPrMqAyKctfQH1Rg
KSCArExR/zddYjFLtysz5UNQFOJwmPtqF5VLzAha1sTQCXReXqzcbH856lUzVTHvfH76hP8UtzJN
kKsZbMy3SMmgVdQZSVIxv8ElsQoEN2Hjsjm3HIh3t/kc7F1QAlgO+6/3uMBkJY2wUQzXMp8iZpmb
jLEYILpluCCfAh4vw5M7zHuAR0lc2+/lM26rAGxB6fDjFtAqmIlx+QX+rL80ZnGbjITNfrSAUe9w
xWYxL+G22Q8g1gApGvsTZSg3hVvZnr5sixl3oG8DIFjz5R4/BydvxbN9dBpqulXAhJ/kthu0jkE/
srJ2wBYqU4ntQAWq+ZoxE/63u4LPV/lgLSRs+T72YBVS/ZJo/zFuDZNWG3BSmBQvmljquDcIYZa0
JWYg55g8gA3z8TBGSS4XD2sYE9c+x4Or66M2qR/zk+RUN/TugJvayqjjtXhlp9rvFXa9Zo4D4uIL
1OT4srGnLCaJZwmdFOXEpWttFmOISz66dBPQiKvU60sB4CKZySG9cMEJvxmNqnhjch+rQhYyaw9G
osP+2wknJ1xne/pVUMNWc0k2cRu4Ku7+E8Ln5s3VyUAmF+wFGvwVPx081idj++CQ/VXTZXl1RLSk
MuIVI6vpwwrNgkIVw1UBV1UOp9B5KkC7MexCDmjrVVY1lTSzi7jhShi1iwLFTBNYlwZri+aiCMK/
4R5hDTA3e3urX/lfdkHoi1xqu40PLIekFw2cOjGAuaZeJzeq/l6qmiqw/ZClUzBLkA6VzfHYVaR0
uQ1e4ng+G9ozrahbCX7/DIgrNzfXhYTZXy3eZtVKsI8ggPcOTldscekXM1ZTMXcYj872pPpKROCH
rFD/w0SyEvepp9T4PkXFUKV6nPyGjZjhQaRbQx9GM2uwHqdu8C85zanrmLjYVdyVZ/NzHWBvyuQo
Ifc5aPlF+GbQ1pq6PucjPGm8RK2C2CPb3lwaOkS4zyLWN8bycTwHhc/qC97GBgOYIKYI34FPmOPS
RxU10agrM3znz4+1NE4l+WAMOVHxcYd9KTihsdoO5aE8B56jhNKoZArYylS6+jptu2x+iM6+uzp/
ydU82+xKXM5A1W4fNN90GmVQKcyORXAc08f/W1WluentStQVcU49tworSr1jfp5ftcDaIVa+B3m+
S2Nc+pF9XTYLlhSeowJigHvW+tRlcFAgKE473XydDNrK0h3bvvbmyVT/uNt+mSCoUsww3tzH4qfR
1d0awNqGJcvUbRE4pnAq9arjLYQwOUdaJD+64TyavPY4GnjNflGCFC6V1tSV4VZiJ9vxNI4vxpAs
3N+6Io9ZWtMovP77gXbwQtzOtM/25OHxAkMgMBElc1l+765JGKnQ5an1QfnpEL93b9kJal72+S9B
djyOCju8Idxtyr0KxcC1Uu54AgW0s0Xncj89KasHpJnHHHzTFk29Q0Vc1ZB8kcAAIw6+jsV5UIF8
+VZaA5CY36ulxNgAjiervr0gMWCRm4YJ3SphqRnuVgNFHy5viFZ1Ru6GtJSA8XX5IJ5i+V0ljbLJ
mz1LPZo2dDfPidoDPYvMgjjQoj0MNx2/FD5liwWfRH3I6e8hFBsj9j+sdjOu9axBVpwoPU+9aChK
hqQyCfybRhfa9HufYDhsPbKfJk/q1Unj2fBJ/qNu98lLk9BFgs6krszqltTMQAyMxCFMORpkldoB
wrVXbIxgdWQGMgMvChC/NmNwpcqTFTYS0+NkPzbd4kNxUiYa1dXYONF5mwBROTwHAJzzhqrq1qKP
kIQbusr53WFQ1w7gVENBPk5pKsPKKr5OuN19Ve+f2AuzrLWnDpYp4AkVf/Z555MF+w0p79GJDGUM
cWNx8DVMFBgvTLrFAdtUT02XJoic6jZMYrj0HdNrv5an7zyAIJ6ogV2LuRm0I4+N6OElt/ew/SN/
fIRLv813KnSvRghsjM8VFsJUP80WnluxLL3XAguRRWa8udpoo7fYV5DVTJ89nw2GYw2nM/0aUjmr
8I0LpnmUdXPE15jRBuf2OTHswAFcKCp1ZIYLL6hsFUw8wout86Gi8dZCmMicp9GeIzGWxzQFk3+X
wyaXC1aEBkf6/0v2woDdnYomkfdfa7KokS4408LE4iwxQRC/iP6knjHljjkPzOqlCpPyn9zM9SEY
4Mw2hOPc2sbBDO39Tcw0ziGBh8ZiztQdzlSI97OSG2pwNU8KqYZ4ufdvDG4qIB+tWheUoJHOJzK3
xoQbYBKJGf9nXONJSwwuOp82OgmKor5Rz70Ix3H8gFAnJr+l8YcC+MVgylGLHoaxQF08hxpN2/ML
3c4zwQSmMHOSAnmEm7xqZmJK5cPBtVoClbUAAEK+cAQBWEf3QJXJGRiHu8jVIm8xqaEamy6B/KZX
jqSckXQWs8lvJy/z236Fq743loFKGbgPLNyPjTl4b56qoIvpXrL0nlwGilEL8pX+TLSMGs+IOkX4
NtZUCxg8aXIHnl8UzPrfr33C1BwPf1RoFu4s+YPPITNClIABxvqrIMP7iLiwqSGeL8qFNci0LgWt
nA5EGjWUQKCf1Xvw+RfatpW4CdA7/7WQ+O0a2VAkR/AGQuteXZBsmPaMmIfriN0GPqtEcV2akdnE
uXZB/tLhI0imHRBKCmneh4ZQNt+QT78O0NKZsixjFVbuiVZSNF3R5++k7uGrXHDA36mBmU+RcvWK
o2F8YH9HqW+1Uyx1EpVi+r7GocZzhnnS3IXFIHe21+S7iOGcm9ulueiP/UzrV8fqEIL3F+8P++AI
9iJHb66ejKPRPtA5J11q9P8udR4BpAxgx04i26NH6WSIH1gd7pOcapD1hB0OVrVcXTNXzvE6FD+U
7rzJf7ToTBvXORdg2TW92h9hM9x2uWkFUBSD22GgbLgjwXRMpt0LZ93MMmHKCUAHf9fp9WdStWgz
uYp+HMStrdm7FOq1L66WOkNz/n6ZKNdutXfiTQPetBnnQAd+IulhVNHnZ4NP+LY7jU3x9Lixeu2m
86IHOIYc3lb1lhmAUAsZTqW5F8B06IcFmP5trArtvPvCFsf+0ytryjT5HDHlRJWZ4lvjJDW0o/Q3
DKUqbOxxbzX9pmVaSSveFBE1wcb00/xG+9ELJ7VIrHqF/vc1DHYKbr1hiLvlR1/bthqza8njqqvX
veVOddsz784c9FLH3KztHLiY8G/DCIP/hZcH6JPTeUOWLOLjGeMvHBUi9W56JQcMQVocvfb0hFNf
ncw/+7NjY+NGwcCyGm+zM+q1hyP4DrTbqMWMMfb4V3pocik4ahtZBPK447mD1ugWa2ROZ6x0HiJA
1xmlfmGSGUTI1C+inx+RInkNwSREmwhGi3b/7MvpXcwUmifus9nKYqHX1OmHMP5eLoXFeupulFk0
zIQitMTCiZtyB335Q88pW03rNQXAOQomkOjj8XztgawKPr150uzEwdSrxz54OaVCdBDLD/LRk4O1
oqmoYyP/EdkDZzoxpbuccfNdM2zNcsjVByg6Yiawp9RpqrjTfEXknFr3wlt2Gd+ruJlgJp1dckla
EXFtxfFuPRmRF9VXa9BK4oph0JZYIxxs1o457/ryj5XjFLVOFcbDIJnaJHQdA4spW1cn1NTe46TD
AaZrd4s0v7NOoiI7LK4KKMH7KgysSGqfbrdn7rccvWxDTXBUA7piNRJEUVvZCNtCUhLlS5m8qV1d
AerrsGCyimNZksc/Ddy13JtGFgji830RymfR57WCbsGCqFQ1nWllarLa9s5F74XnxIqv4Y5D9p1u
utBRF/W4jzX0g+L8cPjWAfWp56dWszERKdr1zNVQADRyulvae+/84epX7EiNkD4qymPqTlbkpTxU
yvB978aqOm0HSA69DdaAaXtIvXNdjOTdYuwWoua1bsQseZ61P8xcRG3utpWu3LPcM/+LgDsTAAyQ
3d3UJzijFuDFJV7EukfKkzaQrEzC40kp5NRc1rAbT19II9OZIMtv4NGCuKbo9vVoubkzFhQatO2p
aewkrwM0cORdoTIV60jfo/y7kBJqJ130KJTrcp8QSWSJTT8hB2DwWLMEvm8cesQPXBohAqNyEJDa
ld6aKKf3PIbGSv9lBJaYv7YvkAl/elE4T4D0GCMjcI876mDsdL0gEhOdqkp3z8xZdjKVTSqT1wQp
WbW/CDHFdl+vtZBb01v5p7kCw5ME5fFOFA25M5lUs7yJb/4fU+zxEcCvFsl0I9/D67RWkXsp2P5l
5enL0vst+/Sn1Gnbeyxt7N5IiHqvZN+MAqQJXM28zRc07oYVgm/tish3T6tbNv8ryiPiSrm/Nx4k
mvGgAvrzm0DswLSnEWB7iIb2CU5bDFPYpghZoXq597gE9FpB/ywF9EfnA32S1Pnxp4yZCKAdUspR
Qcnax938T+ucVzztJfT/KjGARVL35kKHCId13qbh1qcDbm4GMwTRvFu4GLd60UJqhEGLr5PHOO78
HgknaRBtYoQ186Aya/ZDjwe27eh0taJRJGqjOuwa1ExbLxZ2pu9eJJga5vIZMFYXCWuQJNSWicMq
8YESdhI6K+5FIldBYvdJ4C/YdaKWZCkMitKooa41nzvYo+eWJ1NRQXt6Zrjmk30+mcPp0W2UgdwG
215lC0bzjDNBVSKy9vWDBmjVbfUfU3JpPUS+5NiQWx5nrS8psDOvXpPLRSbZ3h96UiycDNBiaBX+
b03E02c9E3NuX/suYrKuXMbp0yGok3dMhjtWmEHhMS2mfdJXfXBLkSWgIuaU3wc4RtkN+WmWy7zF
Pr7rsjJa1JjJGUhlP3lBkq6uEaPoXmElFvT1kk9XWPhZLq/fHaDDGCoPcuEEDZgBMNwjAdvuIkHA
6usOcc3QFptHZ521XoSpK3nhn04t3/raZzZA9+Hm0Ixnyq4QQGQzTxVCcyTxZQ+IMEzHIuetAeCU
+2XIlipCaUn1UURT3/N+ovGTwSVAfPN3rJxxMxnZ/hpFOluA/ztW1h6NOoiUtXSTnWq6+TKnfZg1
7tLkXHY5wtpfXcibtP0xcWNCwrSXIoQMQaEirlQ+rhAoY9SqMHRVouyyt9qF4pENKTaWOkYg3PKw
zkmZMtMUTZKNGglFk933JKD7JC0gQycXIiqEpGJjTsG/oOtptSyjISKgnns86DvCmA9RQs3Ppkbu
DMeSjwBhkl4sQSs0gGynY8Ppv3wOzRKBC8st/Jg6my12uHH2gdf2J9bxaJIJCD68zZ6vych5Vexh
Lj/zhdRqvrfJwJoYYAdkmv9wt5kPUXyP54ZM25KaQX0p2U0GC59nG2A8L/1RSoqXxN1HWuz8Usbm
k2HZYuKkLnQRF5cUHxyH9BjwjOkLEpIrMImC95072VCaO1WhEuL4M01XXYvPKzsbbWu69NazNAc7
JGcJ6vZPR21uXwz6ld+2kuxCLJaon2GJji5iWu2ihJtoIuOWdSrB8mPA0iiRyV1+PqdN7ct87efR
l8lwJoKndqR7pIcStWpAdaUefjcFM4duA0J3Wr/fqZ79bKlkbydzvA1nxncWXYwMcL6PXBXZW4gT
4Vhc6M4mByqrPdg8o1uvuuWxbYwgPpDD0NVIiMvbDLyieNgV4jBwWE+mkkCm0pIoPZX3Eh+f37IG
tN4YuC4nMuJk2ZRaLClgt1NkzeL6Sf7hP0NODEO0XexpRqYOeOvMC7n1A63QAgCIhkSWwaVsDKLE
LEuMDKSE/OPj6O2CXOZquKSkHM6LV6YTUeGBnCYM/yeDFCZi2ZllC/WbPivvLn3l/Q3pNeLzgN+e
29pXIZHSrevQCsww4BpaghunwYs6rV8KrQY8Uxsl3TOhIKtp17Enk7zQgB7KBmg6lYIjgIIXkQmZ
6FqDAi36PLFMrvEqILncAJuAuaZ+WtNoIZB+C3Khskwf5SEGpHZl1sGGyukKwzyoi4LkW9SP4FaO
qJ+Oo2wnklnX0j/Fe1GOmCB64wRdHJ5LRuo6UOPaA5teUIRW4+x/7P45Wv0HkYe//M+ybo7PER9A
jRTQFFPwGrbSFc18G8m75WacLuW9uXYGGccyTnoH6wfBs0mnj25VEsgxQP4zyKrhLtC+PLo7BpX8
MIyr8Uj0iiWLm3PUDWr6qm0OehTnHJ5dkIUe2uijVeeicvTkzShpaVs2O8cZ1xOnEvL0Yd+hoij5
RdCAqbgjKy3uo3A5wFIdTs9ZICfuA67d24dR0GwnsjXRJwjOYUk3WOALxWH3tiiu8Iydbwi0AB8c
KQ9HuksH6aBc1+NCgSrkKYSX9UeFrdJxitXAzVl3NUpMNhLfn+/n2TUZC97lOsmGAe2B361XbYOZ
gDzQnvAkFfSVTAakKmPSAmNsdKh7ClHGgiXLoijNP/Mc/15YLmhlj1KqWsfLFs5IWI2PpIRd5YOS
8OtjNKJkmTe1f/Jm+yqxQtg/Lh3PB1fCSlIASQYuYfnHd6l9v36IF4+ellFmYHsUHTpKXNXXPRpW
JUGBBrS4ZKH3ldRJHIaury00dntSkOZrzzt7ATg3DzgVqfquNU6OJPmJ10kaMhzYd2RDoObidFhe
4jFzvImLmxqCopCGlCfBJik3LYVD6AHccR3nD6JdOiMdsXWoI94bSnbPT8bV1efNPjjh2EDWc6Bz
KNEV6K7PDelKnenn9dxUnq0H9H42sZ7UOMKF4ET+6Pev+L0TNXTIqntlWmQjj110MYtvggdsfsU3
RzbCZI/+n1LwaP4UvQQl/SyFMYkKnN84x0ck1HPYJNzo0c/KeYWfopw6gRJ5I1+QV4sNiMe3tUht
kPZgPgYLm81gJ3HHWAqW0br2HQLTRoWRCmIXNq2qEJuLyv5U5+3hxhaUPDFxxhu6xUn7HRPgNM8g
oOBbrMZBObNuIHYcaGvdrafL8KsY/vrn3xN3bebtEnzURCBN6C+yJ0bfYNgarEu7PyUgviypLngs
mOyUIvptUwSWTCPG/fiLlSDy82/jC3xMAYm6L/vVLllghQBzWwJpR/w7C0IT0iBnW4vhEJRC1CFE
GfPTO4mJHYxpbyKg3xj0zUoQ85D/XXgGpIKAbbBU1UHG93lC7VjKe3aasYhNyTE+S+DHKOcivdU0
GK+jqjlNat/tK4tNt+y73k6FkX5WTdY3KwQaAwI5L8Fb6JC9E0SXJUZZu8rKoKRq5R3+nb5+nPMt
Z6I4kfDfUa33uxNsWjyf1/oTu2AnS85ha1DzjuE8q+DyIiAJMknfClA+xprN6MNQsQPZ3rTr4UZL
1gKV4oC27eCyeAqp6BedvhQNAxOBOaZarIR2wbu3PMAaepg8/RQkVK0jNQY+PmRdmYVHazQ6zwys
js6INg2NeBPZ2urdoJ1hpL7aS8PPSKQyCh2lLuzMHIhQdZ1yfe5A0EwccJP0+KD1/XnXiZXcDi1p
qesQRXeiiTu7X1Mx4/kRdYAtpseCpiZRQR6cQY1ajtGDfWg4/fnJ26PzMziAjxsGSUCNdPBM5vl8
JyE31V+vLGd+uxtY0PjIg+ua3QyNOA7iGme8PfKDf4l07Vn8E7M3BEWXZyg4+znNQ9nfj3Fa65cE
KoZP/jpQoP863zKkkOOsOowHlmHN/ZiueRgE1JtSMRmbc4n/6uc+q8RWlGlzREuyMwA7U/TtEwDo
MKUHQybj/VUDxZw5lsdA/uy4CH83r8paCIbZyPMSnVkN9i1GTND8uUGQ6nJs1isg68ioHRgwt2sz
9SoLV0F5EVKbY4I6dh5tPMhltqxK3eGNrM3spVW1HK/KafQg6MtfuyWu6Z2Qpj6BBy2gmGOLVNlg
TdwalyWQ7SPLZC+PH41iUDE9el2WLyPcydUqXKo0FmSUlE33VNkv62vYHNShutIKOz89WaMpd64i
b9Y4+53jeScZkNDpb5tszF5NGPgynZj8ZGE/jnqwSselNNE5nrjsrSaoFbWqGiKNCZRRpkpw7558
0s4JsMjlGvZUR+lvwC5sF9RP19vavYPG6r4OlO51JLWZOogzax8zftfLzJ1Opzf/TcLiyVlvvoxg
E6t0wPbDXTVajdL/v9HUT/pE0tgBvKAvkRR/7JtrE/A2o/wVTLYw3XWSnSZew5fP07GYadFA1STY
qmHND0hmFaLPFBPzwat9O/Ga5DYuWNyW9TSOsgKgnfNWkFpF0xUUEoUoHvIWc/ru/3Y/2vjx1jAg
e6T47R6xAaJJHIdBbnHaAVniV8C5sOpPx14Jab1ChQEmhfzqYhfBPAjmPK5/HqibmqFe86n1cxlI
/vt73YuGo5bCsM1sw4caEtMlNZnVoslPfuY5V0/jtyaN3aa2qlYcX7sOaAdo/WgNCfAxBv2Y4g1N
M7OsoK+YxIVJo2scv9Ga6mp38GlMDT0SmIMdTssBsfmP04OHigTftLjyYBsOFX82Gd2MI33+nWW4
r2QUgcTgnZ5VLz2cEybLHOwqrjX1i/tH8Nh7GnktrPYPXUbsDCQZVMM++KJSTZ0a1niVVZStORa8
48fLa6I7uqXCvXiZ+eIgNNa7GicTS7K11jloM0Ms/dyXr4qf3Vp1foil7pjZx0GX38QCHzTMON2W
4hhXRwrocUeNIMyX9Wmv3RlI+HZIHntoA2p9XwWn9crQNxE0eNw8dbp83D3rZepl3X7DbKDw5bHy
rzrBuvDgUJoGpfpjp/x65C38omsS8o2kMnszWVoE+NqLmEkRwvEXZa1mNNtTca1pDuMd+0vb10vg
ar0l9YKw0uXtnjTag+r0bFcGWVvUJdMkVBhSzpsNo3gmGoJ5AmZd3OUBqrvuZx8DNZ9e9Pce4wxT
6ErccaLAP+RcbKMGupSfvfHThvbJMV2bbUewEtTSC9C6XQ9oFy+vo00OR1JyXfSWp4pdFsXZxxga
Moz3jszZgBr/oZRfJnZeDs6x1qVMA3f8qGvjHDyeg4g3VrTEePwhtpk05BmzNxeSRo88BJt7kWl2
Oth8L+8bPL1oOG+jsWPwtmMHc3RErYQhaQyV59g9IAaAkmlXfr+1Jhr3Rco+t/q7J/zq0QYg5YUQ
JpUUsF6I5GRCWWOJHtfSaJ7RxKv8RWZtn1+BwP4hMlCoIhDBlTGzTy5d8uHQ1hh2aLJu7yPCYXyH
jIhHFEcNRUT0N5tcwXrVg6GGXgMqZRWefF7vgJ5q6RjsFsvVa+AmSij35LJ36XgovvBHvWX291RA
7XEf1zbJ+Mo2aj7Z99Z8CwVhgHbVaa4vNF3US4SMXa337C5u/eajYOyK+ialkiUInSHZJXXfy1GA
jHvgWQfB1257fQFPO4HyKyj+45xga2SGZwJDYzd/S2s4nAT9sCbvEgiJ3sEcqDWe3/8TuprbaSLg
RqWhfg9CInVf8xPkZuYL83qsx/aBavpknxMkPVwDDRyi3FiiVbixHGvS1MVs06ZRNDG67YyNJK/f
PYDz3lMiRFUeTLBwbkRuPBZmsDsU5Tcns7kfPVRxNjMYFR/qKDd+JU/hiRpDUA/wO3WWO2tEebkC
SwisE8Nz8Uaecpa9mvmoVG2PeG1Pu2x7Zfe96htQKwfjZ8emqLFVAHU1fqUHyESPszYMMILGa8R9
SxdIUJREGeBMBykRvyViwf/ZAsgTnjWJzDAldw87bjYwKXMZvLayZNAFjN3Ss4ywCXUx3w0yZFDP
rLLkir+n+e29Cx5Zt8ranqzuUSKNlFvnquDxXjNihfFoywpuRY+Un+OO5qmlP+9+vowj+QkLg/oO
RzM2BQAwvYWq4e7DJ6gJ/sdkB2m9jVqBcgMFAI64ILoFmPxtawj4TZ8VJ/AUWorUSPgilVBvnqs7
awbURqLOYxcS2D0+UvatWDE5K6cmt3tbjFBgRAf/l4DZWEQjmdlVM75BQRftkqmQMU2pz2+YomF2
QhhfMWsHgzPHSZiyDkB+4PD6B6bnZzxJM5jNaWSgPDXfP/GKbF3W4LogFeSLO6NlKdBWTmKLMU2y
d3FSDcrCUK6YF2iV75jPdzN/WphDYCEQ57BvyuBUeDHcVfz9VF4E85l7BTN8f8N/IdDmi54GBrGX
91+VluBVqgM0nKq1/lBNlzZbWgPrZveQEWutImk8kJWM2QYg7tgkdLpvZg9UUAyL6zrHVYPeQTQH
UKms3Prn5jBuTBjauAHOAWoFsvnbyyBaDER93thThLzkCljr+ZPp8p6wwYusuFM/9wyzy5iOc7m3
gGiKqA0UpTyFdFkALU+6riNoy+rJrQmbMhN1MT95HvITdDLMCAwzaN6oKOVW4Z6qTrflayemhqqZ
hlBnvio8kex3f8NA0j/Rl4CZZzzqPqVZojFGHFoGn2rPSbfCN7yaNQT2SDxxPkLELi83grdVPOk9
6xO44uUZQDgZUwxdqNzl/82tMJIiKfxf73GZeYRPyR2DHCNDG4e0rHS8WGfVcHf2Ef9zzVaIMyV1
w7BnO1zOO2Rex5Zait9KAQxXvrKXsyzai6mhAQDdGx/aJ6wrp607z5ZzV2edFykSWxVlmaV0hN1U
bRnd0IeDjghVj1amUCMkMwh+nNxdv82Ki76u7S59jCxkqdyEXdIKUuY0k7BI1il2RYBqPljL2Nno
S0fBjQms7Y+ILI+d+B2qP6eTb9CQUZBHoBjGl2j+/9NtxjZQCtJ0yZeoSLZFae5te0+Q1qQfgBDc
FvHD2+S1aaaSOBQlxs847qzYOBhskXlV1HN0fneUG7l+B4FEk3SvIp0K2G2MFXJBHpIcijWvnRae
zVsOKnmKFmTYmc4ujW5tj3aZEbzdFTMtS5M9CbfyeGeNjJOYeqY5tPakyd2Z76ZvuV/PE6XjS2gw
gdqey1ZzzHzwdDaVCqHjIInMQAsdun5RXGJyN/wuaaIGyaPjU8DZXqnQBpH5w6reznKauWO4mox4
LAjxWuwm1jjlt/GVfZ4vUidQ2vL/xu+WzXL/E7dz2/AZNA68poj473/ZF5d84nF8urbioH52qMmZ
7pDbx585sIHyAFMW63Q4FKw1+UKwj57rE+2hkESet45C8CtXx9IQ3mXuAGHzvZKTHrSvQcR9kpCx
grQP9garts+UocloXqcu6DpeQ4xBboZ8kXDC2WIIn2bzDkrXK95Ls87J8M0Qj4Rzo/EyEGNjqabU
Ho+/H6Vksvpi13H5vIIzm7LWXdAVC5H0d+NfNGvKRow55Y/7C1edd/UM9q3xgEvuACYxnxkfyX5C
yf7LsFblIglNQUGsiEIDLJPF4GB2yGW/HfBk+PLC/gLzVcZpWPC/yn02nY1D2vf2P7EJO8cBt12O
PiZoadNwzrkDPt4dYUFK8I1wUP26HgC6QU8rLuOAddipyyeiH8qoDzrxzARlg5vWl8A1MooNv95v
zG2InVrST5pcJJmv0Yi4sv9mu5CpHGshr53Kib8yDwp349xRKf8um8Zo8QoMVspWj1htRJtpDTBo
6td4FIH5m1iIX+E/UOQL9rqyCzXIaHySc9z5U39lNDILTsphVdpJ0qhqWU9A+0YmRrIqpCQMFEGE
X5AXm2sPKbhpfg0mNX7kNNN6gKZYXOns+czV1J4dsAFUX5+ZS1t4e4BUpRsdUkuz77X8cK56gmWU
53YfYs7RLSzNsLj59O+xun5XGQp1mvH8MLnphWBWiMvCo5Rgugj+zeY4T+uVCYmHaE0M5pltXe+a
qGYYEHRiY7V2ef8fPQJJ0nvi8Zh1in4DuyFtBMsQeQqJmTwJJ6M7mcue3RftyROfTUtLKM66Bgxm
Z7QAE8Ce8ykMtDLB9i7WVV9mf/cXIMSmqTJpEAS6pNZjpH0uCz1/74wBmd5L2cvHa1hhwAVWElEM
ZE+dGJXyLBwErZXysZ9ybd8LPs/vRPbFwiL8ufM3siCrKqcwzjEJokKY5/KjOBngVgStNK6+xPwv
P0W2G6vlp95zn3B4JpffD/L5KKixy6i9lgzKuOJHwVTTmqD5py8kJuuYF6JKknw1Odz7w2yFZUtj
F6OyKhMw47qqjk409kB7h/HJ73fUz8Z2oqwAXijVZ/AknWBgZ3jzUFAy/37bkcz2qbx7BkT6+edY
3kbBOX77El6dpHe9KvWTE4oZNYXOWlJIrn2oEFGlP/gBuI0BZhB3VkdEZw1J47H/0OJC98LUStMk
QKp+L7FZTqplpVHN4u6E6Gsa7Df7sg8mG+bi3eb2FstRIHyrPYmim67IWeOTRJqRhWhY/DfBJI3w
lUE+WvmdTKZq6gVVlQADBvl1YyWpjuH3+0MYJODnc8mB0xSY2Wt3k62lzlFZIDhHm5EFv/0LU745
zOyXek2bPwrabJBhUHoNcRxjs7lcrSLBrVtB9L18f7y9/xZtPM73x/vSw7eSGfuvOIp4yc1UCpPj
h4BaEEi75LrDNHePztroJLbGKl0ODxJ4N5CsUF6OOQRGl3FyMl9CvS7YQnRV5Qih+E86TIeWT69q
bedblFZoXWe5X24ncOVpXr03MsItaSIgcxXS9S51Xo1oeQoqlVfKYn+e5jlCXx5IuBrr/h8rYw7E
uUHuBU+v2ln/ugOFYPBUJ9RPxDJ3pB5HI27CEe580ggF9wX2EiwjiDq5wJ8531EmTAJ+Q6D1PE97
Hv9gTA9lPI2C4adfdT/h9k+uxvaQLYX1gF6E+PflFHATGmH+NK6Ng80a2Jco16gM1ZhGoFt34kH4
cPcj9PRqbXtoVtwmwGSG3KZ3ZDmhFTA6nmcue4pIU7O94Vk0zAeL+ElthH5v+NRKD9s/gldn2lVz
uRD5Mrm7x2z642VJpMfgynfaT3bJ4Ilqe5tdnkkrJzCOBQ6+ZF+uMQMfZG8eGbyX/8vwueUVvy0Y
zQjRxF8+tU357tlXXwXZb5khUc3srPhpLae+a/Kn9rVnwsx29g6akl1npbn+7/Uhfs3d0hrWina1
VB2wvts0t8e70naG8k8OrJSIaccTr+FuIjjoI+3+fzoaF62rBcJ0N1Ddqk3mijcWk/i+Z5Xc6eZi
JCtmFCiZlGUciGzfjXuuL6AyaiJTRC/D1lBNGLl/6YcoB0SSo49i7aFL0bnd/s7u973oFNeGCx9T
q0X2sYSBD/3G5SpHAF1+0jkZQ3UHcDK1BzPJgZw42RzbddOsS+vAPXIAhaluvtJY5D4wPpXJQlri
TWRDYKyPERyXBGdAiw7PazUw1Uhc7hdJSIM93ibMETpkcKXyKSWvsS7nA+nkwWnNGVX/oLbwByo2
EVgUsVDyiZZ6poA49BzLjwWwmUD/4lWTY8m9klELBlM4HOlE8fQYuTWNimik2ZoBFXsf3MXgXWN0
9Br415NhvWT7QKFuVTXZmoZ8pg93WskVxKJM3QrMTKpAp2DU07M9UXQKhBsKUH7MHejidLtIgbyN
i7VB0LvUkF8p/ML9mOoUWNPR33BMqh559CNDdFbwxVSUBYapyQhpQ+VLyVis2Q4JjVEmN0EfwGLZ
0QUuHuAganmrZsqdz7PvWZfXhpe2dCtmkGLcB8GtRisl6Aa6Iu1fcRIUsryymAErsQT5fFCNcMmG
b1iNlOjfqKZ8SfNkiP6MWrAknbrcLeE6/Lkr7VXj/2zUi1YpyaLhwYhQ63vPHiJtYdPmZZLaRz/C
ZNhEoUWcFgcSMGWjAc+wiABe7/Wq9O0w1Koj/Or2VtWzidR7Tnaz4M9HKGGirJTlp2fPK/9VG+RI
a526s/jav6ZFsiwuhs0qQB58G5C4Z5RbGCaShPUTAVZ0W3Ad1s3K8bOzSMJ0MCr/hb/hRrkdrLGT
VXgrkGs4x4i+wQlCCwdDIAk99ha+IMfyhAmWOS5R4iL/1yFy2e2iORccEuOYwT96jRD5M0LoBJgH
Iwt3hHRjR5sUsVXMdOlC0GbJMlSwvQmaU4+LOUrmlxDdI+shr4Sdv8FVg3hsA4PjSzg3RLAyUs8t
wUWZgEB3UNJL7w9BspY8vKx3sA67udHCDFGdwVf4BAnTZPQR08UBggnPZH4OHXHA8RzwW6v/5c73
1krvL49Egv7aIKNgSTfq53V7xCaiP4srsxrrG+HPTOe5aYvXanOi807p/AEoSadHpNrxv6zKDTZB
WczKJKSV2Fcmj8j3GHu6Vga28F7k0/hLUb1BYdrB/kqegWaan2WmSJ8QctEk21RO89+UDZUe/B78
F9pYMDOeFKK17R64Da3vyh6YxQ6+QslnBh/2KtbeEhCD7f/eOOD12fJiM8/yO7qJgePX8dkSGeFF
suSDW10Ph3pOFv9RYreR3yrifXrwCFZ8rGbqQScqozNTUEj7eZIJU255RC6UGBUlBUDgfQrdU2+n
wWGH/xxj2mPTlCunO9T9FYnHToSGHNEKWeOJtJ6B27NkMVGd81XzWKhHOM5VtUZBsX4u6WCiwUPF
1aHICXQ0gWLaE7CsciEVMxzjoMHkjScV3wtxlcOGMaiaCeMuK8YZL216K3luDXru5YEMrWr24VeN
bxvSylWfpDJvNoUUTpXQ70D8+BMxq+kkigRvO0enOZEAXmYzCH8Lq7pTXrXVdbKNPTJavrkI8+Dz
JztV1mB0h77IIk9coilBOepSeRyOB4Yb1Ger6V4c3MHMe0wwZVmEl9X+kENjSJ5zGsAVh47vnt0m
B53LPXQlnfFtZeCrGc/a3Xh+6F9nEDdXlyzML9+osz6Pnw6eERhaKRfnF5XZ6Bazq9U1Zwhyfs7r
28pPwgQGfTBNPdKAEiszBd4wqXsav5nYuYabAvI8AtUkkieysWx6ZU3Rfmb9XwlHTJKcoUF27n3l
Du6DIvlSqtdweJ+dGNKhfwXP5cbouxgpvqU6CoALecTmHq4RUGhHwHAzkPvzXINywfw62A4g/5Og
l7yXqb0qB4IiaugitQSbgA6AVFrMd04bgLzKYK9WCCoY88iPKjx713ZnfSv213iZIgMxLQIn3H8O
l50kr+x6vVG6CusA7/bLdeW7pDF+UEdlAVJnVz5JEb90rELZjLE7N83zShTcD6+BkqJb2lNAjA/2
5r14qe4oK05rHmLdQ/IqMICLSdxmosH+REwu0E96aMF1mK9v2c5GS2p7/LFJWHDjs/LVMH2kkLhb
n+NbosariyyNX28GglrfjtpaJPQv6Kc3xhH8A5TNxs5W8XrRCiVi/8S5pxP0snpkK9ne2u4LAiFd
ACBHfg0Q/7dnBGd4ErOBaixjhnt63m9KEw5DoWQVBnNiuoWYpyR+Y+fYW5gOugmBb8MmyI0okmYd
AozOdoczBYXhzmcBCHQnQATqU2YDkT5Mnf/+E/M+BZTmVs2MFj5subGBejK3mntQj5tT0CEM2niP
Ie4g534+se4dPhzfL7B1D65L3S/DL54XPsq45rJ+lQGiWYqrf/4r5eterN8COLm32YGeMbCon3gw
/k4KSL6EBXkaZgATpXhAtybwu06jwn0RuEB+gVSesHeBBRe+Syh+uBT1037fjUSV5Z0/e5vaTMfX
VzrW5/0pNetDgcr9ajz2NrEv3HoiqoA3T91MRsF2swE8qi9cxwb+AtQc/v5Vxn4ku96kiY9rT0Jc
kKJS1OeFVV1fd0RpLOLz2eFfRqb2v0GHYKTaCRCAJczeR3XHtF6Fa3FDPYZ8wXBVnJv081AZQVZh
L5pE2WyED6rU9I2QKKtX/mIGG0I3VxnsBa6UzLVLTDSqLKi/vExloQfLU4UpJAgMhscMfsEHmV9z
AXlL2whsKMBNIw3keWSKmVo6M7YKFQKyiEVfodMDq1pF02M25QPuld7bQa45N0Bp9G/6y0jtOv/2
dV75BDncjTIzQZbAA8gdsyF3BJjnUbO8ftHlqSrJVS1/8bxRGjjdgT4Pbwl0HkL4Hfc9NdvQiv6U
nwb3+WL+4aoWNZ2CSSP6pEJrJQG4o9493Xl69orSzLqfVxpVRpu2YnWsZLVV62xVkXfdUA05UQw8
40BSz6oHimWRbXdy8PbQH1TJy7L3pyN6xCCBF0UaFiB21GzdUjxmU8XQdSVOTCQYBGWD3FsyvdPH
voduoMXGo5s/9CLGbfZI151AaGXGJ2yzuydOtLQ6LMQ0/UWfFWxn0c2IkFi/eYBhY28NZvAV3hFP
5AY6YC6XhCz0Qd/vPxvLNnWQJtFpv5DKySjn6ssYWyg4I33JQAy5AfOy/3MeIm/uK1ZclE1TCPEX
y5KVLYMVuVAb9p0kXDFqYwDCbXT53fTggI+0re+cz6KDncLoMFwqfPBBwD/u0V3vh5ZLig/mim9R
NUiDxctrW9haVj8BvNUbvmGwRx2P/vXcUZjJh825NL/nxqaGTWjzgsNx6LbC+2Vs/hEgNwnbUQeK
8rj0FuS3VUMpYqv8n1E7TzglxsPl5bMLEk3xGGJmT77yRbB21HcLKuy6Jfm+iQciZ1oOsz3vqf4E
zTMKeRE+KykPOafKKl/w3rp841lsRo+c7k7bWA9L7/DfTpJhgQTAXumN2iR8qoRicVedt5XKLowH
VjEez/91pYLBjBTmJKig67pYeqkuFTvKgJ5v6bwchDe4HbYd9qEElfQoOaIm23DzOr/jCsP0fA1b
AKyOYPOSXmWLFz3OXpop0XsSuFnqvd6qvu8k3fvO8TRkMXKDUMf9APAVGNE8qyvk0ctprvCWDDKH
QYvH81VXFn+MQawAqU5mPqmuhPn8ssdJMUWz/Z7nL5/KyLYbSCSgDrINNKcVgafDV36gNRMj58h4
H3TQJC0HtwmDROmjJfSTmvjJBbsNDq19MWf+SiVFqZpTB/Mi2TGGT8fboK6XLZ2ls1Kv9w1DFeer
2o8Qf4hLeQKvVAWGw3+paMkpfAlbTEnVOWaZX1fNfU69Xd2PyzpgVmhQr6Z6X7KiiZB9Y+/yuTJR
KH4A1Wr8QDodhkQ5F2X3rNageAajWEBIkmOaS+Y7VpOCQz5NTPDak9dYOojYlzbgC67n8eifb8uI
gdk9qR1H7rNAhSkXDS58LL+D+h/GKhu7mkSUw7ggMlIn3CB/xYq4u6LV2k3Y8/QQAUnSuc+BVWV+
EYlWYKAYBQQy/84RPbJsIlqCua9ExceFCu5m+1Fah+7b2EwYHMqWzAsZkO741/iHtD8fBEEKwmhg
z7EXBeuZRXgFUYiG/9X+kxTLVkA3Jf98feMJXpXK9C04CNsCFXj9ma9mfVUmSjM40rsudGEqEEBB
Kd2OL2xLE4ZmjI+gRiLvxyollylTHONBQTJXO/Ynqjy7NRv+pWtpxDZqiTqFubuV8V+UEU8Ii3Z6
tvm6hHhRdL9tnWIDkxTITfY2kXNyBNAl/RmermGu7n952OgVl80qLY4w93KHeRMqyLIg/eBVzOUq
Qr5Wveopa6zzLms502WMzdZN7RvHhK2u6eXM6+4pA+SVh+5Bpm50qrLXkgOKBV8QdZakhaihpIY7
U6/D/nxH4u7nwArGTBOnqzZURqFc2lCPXrm8JLvIpE1g+BSuTTMdEwK5QL/MYrhxLUcuay0YKh9m
1zyWLcWKgXSL1hC0vYTJJ3i//ctRFI1mLcFuVcrn6GbV1Eo2xPieFsvIT8UyrfAAUijeRcJV/J/E
LrLCHwSSuSNC59jvyP1lEydwXztOpDJuni3v56WRkt1wO5LzJSM/rkQkABCrwDfSelu8Pd/Htcvy
FV0DDrWPod1sdzr7fwPr1cMpygSiX+CUs+cdEEwzlmbY9DURDM1JO2WbYEPyXaN4Zce/aKHLQz4Q
czyYXcMVRC8for3sMvZxPtInaoZPg1ZIX0cVpNEr9a8dqQZZph03bpWYDbZtKwEBHWYUCKMB2+Gi
HdvzmnaSIFdW5qd9n4KtUITRlXOpH8674REIFFjxrDRMzkHgQtezumGWGiz1WWO3bmvhXE9zBlXV
IzweAlI415/eYAZ1pxPTZ6mz6lt8LPD1P2Uyoi8dPB88lWiNW8+sqCerdZtDGjNCruCUbHGU80T7
HKVXZ406TUXx2O/CPrCA1kPjAcffYsWvahZctvZ7w7c49lBI1y38glmoqVCsX+3nHfqd0GoS3kCr
UriBVGemlrQj3DueLI0B1l1WIQtUqWAIGdGjeXPbOMEMkJPyAG++jy0bvQtyFMv5ewCtYXzqdWGn
G50a+YGaLM3zS4Jp2qBMX4uVIdfqgVHVvpDu8E3XOuWwSYopZjtoqhJzln+avvyc2rZUAL8lIc5M
7k65J8DuMQhOOxUp+UCszO6SkNZfTS3h1rQgFkRJQK2PGo+iQV38naGPlgjGa1hUR8r88m/yj/0z
z/cP9jgM+4TZT/QBdsDhiZYuKTvf7sikpqJ5Jgx6ywLPgZShI1y3e287xzPqXjMmBlwogJWJnsoc
OK/V+jvN4tKNCTAiFndOim8Scm2HiPsI8a4az2OfVS/OucohWj6br96+YLpp4d5DyGdam/sGFfFp
0KC0rJCTqj1ZttXUKVXVVCxHWIVmMPXylbxuVOtQlqcn5Te7/H+okOBV8Ba1onSoEwduTPElHHIf
dYbvVuxzhJ7vHV92zTuorAR0uv1WnryHCOANOXUx3dFrr2nX9Z8EnRF09jwQC9+Lpxg/XUzvEfDj
Jp7nhhICvTnSFcrqhEoWNto6D12mMMydsb14AJVbJcoEFHAby7/wWOJ5KQfIMhcQqGaqvf2OeWUR
MDLEfChOYONMQFyHSJfijOdSLuOgXOXmZJZ3Yp4H16GQjeJQvqpAYT6fZPOAsMwTiiXGc8la5V+4
ZslHqg9MVgmk8Vcc26a2CKoLBcUQsM6RkSNn503Z5jh551SZGOtvveJ2x7TBBD+hg8Uu/CCyCC9Z
2hvPOeXaKN3tOZ0fPy/NoF8MBieheJOxsOTsB8Yqcsuz+s+vV38m0msridZKpMpHGupaoxDPMRGj
VHy2IsSCPmW4iNsP1K4Odt3JAeyg0KU08z7gjoJpX4yJL1OaW60DZCNKVFrhL8kPNgbdgOPdEl9f
vNLmGq+JmsGu/6TBfvQonhpK7z/mlIzZrV5hQF5Iy55HKFU0M07FnA0XD1zcoAiJqOJtZuEJJSIE
V0vGbBVcEfRiDdaEUh4+VrVJ8PpnfhUcOEWBpgp0gvRANzxCYV6EqfzG/KWukRVgj3dRD6ZKCSVw
ChplQ4UVz4YS0QfwjxTMUMl/cTXvFtufcINlQ5n7HKBXD0EkDAF7oPAKj/XbzFGk5GbY03faKAEE
4nAm0p0Le69uU4jvP5Bxq8z4KsBrv2XUsCVZLvs/BY71jX/istW0xhelgKFkBk1OjXROnBuSC5Qo
GeJ+4Jd9P6ePLKBAc1iQQQG6G5BxqeLald7L/CQsORTqIG6MgUTw4o7XjPQoHtpJMdmdjVucqieY
akqmNlS/caA1aWL+mR/CEvsUWAN8sC6ObP31BUxgRDc4Zytivi0IUdUeOlw69QbjomgqW3zVZmsm
5XZnJFHniEQ8oAQrTYvmshvwry1+JBAeCRQi66ONY9wMW8zHiIo0bTPESpb1rgLzH+nMqV46usjB
VH+o7hTUNwQ1CHBDQ7pb4frOCVJSoGAELtIRO5V25ivbJBbma7ngIdO030x3SW/2UHsKXog4VMxr
+5jdDFFL181viGz1VzgCc+O2Q+3ZXzAWXp+5Sn0bGtRsS70srTK1Z6LI7Hw4/OdE1fNDuOt4Iifv
8SQNn0x+uICt8dI2tgekh9m6UfdNdL/kXapmYQ2Zp3zRvviEe9ifc8RWhVsJhcndTROmGA5//9Mg
QtYpPyD7bFND6q64P+sDtnQFL7I3ZImqtfo6urI0LBwVs6IZy4Sa+68wDjGDeM5iT+bOijt0vrJk
CeDvGT+c/1KGUK+ejRC0HkDXYaWgOpegSHzQkXqOi+lcg/A2m9M62aaqHKiWZ3u5Mmz2e9JECLZt
oOgstty15GoE1MIvAKt6r3Z3cifhI7etRfQDhtPwOm1D75fhreTVVlY+klDjtRnDJfezR3zIENbv
4QR4YgONUgf8CTPVYAQP/18vjGgpkLeQfko6bSk+iGI6Vf12LDmiK7wTN/53im8fUu/Go0FUJpa3
UPgErmytxdexDDDQ0X2jY1zb5KoQEnW37FuLP6x1J/owGRY+c9FeAORlz7Djv5e6B81A+NGu9TLd
8+F9w2BUdGZ70mQe9zD935nE7tg9rgRXC0PcjMBahymf1YTYsTxCTrV3z76yEeTYukAt58Wnd2YN
M/8onR/A40qTuzM0MtHrd9V4BT3Y5FIv0rfkxsIDHRvnswoDf9thqd6BeGeH6jNaL1T1BFwio/ul
6S+DuzqJuDGCP9vBSWV5DOEGEnqdlCX9TbWSSTnYn3PA/3AZg0OhZsFBEANnHl0k1dkKxCkWnkzW
prl3qewC3KPTPwAaEMyZlyqZXRctpSm2b318PmEkQSvQXxCHXBDA907e1mClwGYbVf4eszlsWyxI
xODFCVvmQmk64ERSfWsdhKZTQx8ofPZz52oK8khMBSTmpaR0oLie+SUuvVDOx3d3JpSbdQRSvjoi
svNHkQfOl7cvUHfIsVjlZO7wRKMtt3KEdmC03MnCVBPKXoe9vEKLgmxMQd0WCuVqtmcjS8DUhvzP
a1Sw9l8FY5UUpYZEI6eiOBCVJ6Lf2HJKoyPLFP+2hBm7HeN76fybZE8vurRhHLSio32z0hZrHKWx
L5Caukp7WW/dEjzqFclyxhzUv15CIC+XyXvbOFPxlr+iwxDhcP24jAoCRUw41+S+dlIErmzL7qFp
8CUO7L3R5ah0/a8z9Q7kj4jMU/rIyzN7Tfcjjw+tP/YPUnGC3MjXRhcOaG08S/qmIRcF5ROcuS/G
PilsAeexkICqJ6TwM6lVGWe9tIG4A547BgApiD7Slpq0RATXNzLkqTQ1HspKUHm8/jn/Kc0orfMG
W3BLc+JGxdU8Xk/xdEhF76ttBmCFNoxVGgp5R4OD/qG+i4dCggOUyJ2vwn2/1j+5K/T4jqvV9e2d
SpvZgJ/RqC2iW8jtPxeT9cQB2aGo4D2iz2Jis006Q4kppuYsJcPrr4gGavqDVMzbO6Blj5Ral3mQ
scOzNP56WyLyjVQYIcWk2I8sD4Ks3OApD5fTbRKCJw1MVlIuO6BJEEC8s3/aZq0u9qT3Zf2D3p7i
qvGZXgYgzLjJzv+4NmDLGIq4SnwnCp6HSpiy6iDgqOj0cCZY28kHtV7tj46C5z7ypwFddeMRtE8T
sObx9Jpqd4c2NGW9lCV6w/MO1syAVpebkLCcmJnKL8QlnzlWdyM8/1Ub/+VpFUcMjPuJ5f99om1v
cXCBloDjV28MqiC9Yw/BSN4/knKrc3fDa9r5FTRWyFWodOJ2qtJMoDIGBkvHPemT/ltucTN2uLbn
M/AqRDmIEIf5qqSQXWt8M3cpJH+M4d9+MIKW92mufgf0lnW07SocQ26kgsGwS/AOqSdZ0LW708mF
SGcka8KVp1eZJ17KwCnCJW5i35ipyCvv2G+Jk2drawwMlLDcQZnAWxaPnt2rG8Fx7aMQ+Fhkwtqh
mx3PI8YXErCqVZ9xtCVhtIz9TW+yhPrw2YLcULrhwk7/xq6wsiQ3NPOEMdcosEYW7mpDaARBo12l
hWTK3sOVcUjEH74hqVUdwME1u2q4QGLp7Juxw57R/5bvXE+8H+gLA34dvgX0q2zCJJ96lPvsFX6z
KZGjprvRdRbgbVyDxyj48fyVmDFkceyMJiPUt6tNyZY+h9Rtj+kTEcNIe+yIj7L8ldBXSR2C4mLv
x9AU4WITPHzGNpov4nd179vVqKPbBvNwQd8T4MlAoUdNAKcy1YSGqT94nOq8Rg3xvo5TjuGtWCXd
sseDzmlXcHqTkjChcaEw96GTGPVMdLFecdhZ4LcSp9QgEaxVnIqdhCEz+o1feN8wI+0tIVrjviQN
Bvna9nm4v1s/vZJKu+tX/MDddbhduBN6r4pQL4PzeBIap18L6VBbyXNSx4ERWT/YsaZNWzNSrobh
N9M65Oi/5u5THgSKFUC6x8ztLECs0LuzKs1fHh8aRTr6sJDquXbvWKvbotD18CudKIokbGceleJZ
G3Qr9Y336EnXaaNVM1OfZTXxdXYjAmxI2jbCxkUbiQ/xYxBJo2IDb6bcLB+iQO3opBAedjF1OZdp
DqDJgU5cOuS2cobkaP6sMskWo8EKXdzHvXAzSupEJfUjbGQY9/0OsD9RNInJ/zVKW0XTTlAsnmg4
XtM3mldYWbEBSOOWDKagfkVcOo4znc6SWsQzSjqR+9rjTENB5c7AMDJiQ2nyWkIK6eRr83irbK8b
n9Ehn6YmLbuapeMjWm29rAALLdKO6/XTw2025BUhB/KDBLfiNxwaDByPQsiLtIhkb10Wi0p9OLPd
/u/WsoiSVhqckav/Ev6aZcXHtOynPqgUH5QnHKPzbceujgk4WWmwqM8j+0/0amt9UKlZljALwquv
fqe+YYq/d2IA4obRFi3K06rm2blGtfRAw9Jl18gx4sI9NR2scORvPs1RMhclGJhQY79vInjsBdak
u6YiEcXfbWEuTIGMiX9jNhmNkmqsr1OY3UN5nPsPg26XBzGl8GdL9Mmw2/k/4mhiLpmACYEhOE5W
y9DcvLfv7DzM2WM5fa072bzA5xYM7rQ6QH8IfR4XXa+4N8Nb9ATwZKIfmyGPDs9lMBpk8Dw2etRS
53pbIS7xHa1q/L+LIZZEEO4dzNmJEh2pcShqMLbJU6XNJLA8hKDivmgtUdcVi0TnpuQiyQJpvRmY
yDdhXTKRrSAWrhqxOOvZTtY/hH6JR45YDzMc/06xsHW4PzhGO8XaiQGyr95xRzNgwxNnCfrL5ukv
3BvfANat3WyWI2UidCjmdZNqbIFAUvcJJC+5Vw+PV5CNWjeuhr1hLmvXGFEP2pwKuJ/7JgxudQJF
onfQ0AndTOVeGcTjyGAhHwMqtEXLPPSXJPxKbWLMktAL6ZlP3itCgGHBSrZJ2A0VJzlo6xc0Mb+O
XEohO/fWn9ShwAJrOejKQylRmMWQG+JjDaF+7VCWppG1u2iaqYu+ZVLVps5t2nEEpu4uJK8Ejh80
DDa66QibQZAOEloTSnY/Wez/tL41UR2E37Yhy8lYVC0dX7EIBUXdv3pBoxXV8PvWrc07b9HztI4x
HwyxcIHW57ay4FA/eLz2KGvWXGMUbCPALWU+TKNcg4zHgnxIb7LRoa4nBahnymuRydjrEh+QF6+a
YgTWV3hveunnFAx6plBgjKTmSXPrLBTOiVV9kNaTUDKubG7FHNyP/136jZTsveiJInNyEtugHqpq
3mAcPodhrMp2F9lQeeMVwbE2usaJGZK8i2FECPt3hT3cjwL/OhhniwDvCYUKhpNvLbeHSki00xp2
6tJd/DhqO8uOWSQwcR6tYsn7oc9bF6Nh/6OwC+Ze9rD1BpHX71Bo1ZPOzh2hteHp1gYI5+j0yxP5
qIMEh5by1SgQs6B6qsA5FqEXci64t63Hl2tTS3l2bH203pZs/MB9mxMBL+hWKMx6BgfR2T9SJPCf
UgRY/21azxZVulDOs6wrpYFN94kCWAT0qKrrdgHRMZRKjcup5ad+G1dKV1cTMr8Zwpl+LrYUUc39
dvFcOA0CLznR3TgWZpQWHsG0NtM7ppNw1px0+yRgJhSKrzDai9Ye442GHRYOGl0TA26MMAmLqcF/
NiRff1kUt8aAVZr4QNMINcq4H9eS01OsqdrIXfW4LOXVH4Kcm65si8XEfyygB5scx/D0BvtuiqKI
xPGcCgIZ72DiYajnqRqrAkY43XwdOSHbrlSkmUxujHgAi8P+7h4bvnmr6NeHvlNaQmpX8//y4AO8
HPILb0G2jZCt8g0VpkNqu3GBbZQJfaSHqTHnKAKBPKRPAv6uema4DSEKPFnYn/Z7MFNhZy3SrFtO
k+/I6cYMwC4QyZqtGdflu9A/YcRxwpLbeEbyEY0ADcnTpY0dbHZZBLGcgppv+Ejaq++xbVwMCMRE
DaudfS69IcAaa8n6cjrBgKfCR9JisMbY2XQ52/KRgIplJVgpbflqoGm7PfKiYW8yw1RRD27VOMwD
q1sllu2UVG61nCNaLe0yEd5+ptunO61+ZkQqL5xgMboOx6z+m4g9hxZiLMOo1NRPCL6x0s75bwSe
6C/ESUUDVIYWEPrj0ILBsT0Q1EoVBWULCjt0rrKNE3UgFTsaSiKIcX8LTjcxVD/XRPw2G1kzDZBl
G6nN19/Mtwr45fwyYoIC/pyU9xJzYPJEf+jHec6UUJoTyyQsuG4qRH7FXgjOll4HX1tpvrFp91tp
GWee0DpvV0bucww5KEzk0/O4AJ04QM+sqyxVqLOPnPgnSq+8sBo3xlxhH2KKWmyXFFdXwTH4x0rQ
kmj7OoDzHZDNhdPnLWqTwmZhoUFtJa5qt/7Sghaqj+z+gmwCMERbs3VhxKEkhhQZw6TD+zgoYYWT
SdcLGRT3KJn2BEv6ApuxwyVR1e3/BIae+wPHp9SuEsg/qcVhNnudOUyDpD98MzBURCs2R5tg9n+i
tfsF1hpVRdb59Kh2+AmQhRLLj/yIgKTgKDWk+6E4a+IlgBwhc76aHosRYWsXFKI0/roC6dfVT5+n
7W4UDQXap+btIUgLwbftkPzHMXqF3Lyn4hEpbuJYNJCn99qL20BvzOuUgw5iJ8/N4NO2UCjCxnIW
5QJkZVXHImcFcQKtGHjwgOvGUPSpeczugsPN9UV0E+aOqO7L3yeheRP/6pjXOHSUKtNDPfIzLpR7
jp/be/7IB8ThXsxgg1gzyXwXwqJ9RVXoscd6s/0frVFD/BAtt5o0VI3NWJgG4eVyIJR3/IjVU2tP
qkggHkyQ+zyWOahFho07bgiWN2ToPHfCSTrRFDwUTBXPoktqL4sXyMPWa8NFzMQYOqqQi2an+bMb
49znfuEqSs/4OrfpMhvNUHDGh3xkYP+lnxwTDTYPGWIpJCiZKH8aVq2bTAFG4nLpJf33cvWO9POZ
VV7PIF+oopE6y/BkGc0seBdBzIUEyZZc3trWPLGK0ZvXra10QP+YB8p43ngXP/LjAIEelWcaKYbd
VeCSQ0ezCdSkrRGu3YD0ZovG9yB3cS8yx6AsfQv45sheelh8ulcQ518NqXDtnbwwtzlCuYRnAVvR
0PkJy0aOo+ZFYeeNR9ExGUfV/dasJmSkCZC+2l6ECfI6zvtGn1MuuOP/Hst84l5k9MwBLzdPAAeH
xRzCHGsrf2eFsETPKS7pZ+Sj0MnM5N0Cy1TvYZ2fUykqhKAq90GDP9x/qdRpKdFN5qs/PsDX2f+d
JnBcr9cH3hAN0craQL8BJXYn/a3ycfU8ez/2Yf6zXL3z21XyA8PTTHzPPpeSfSTbyb2Wqvwqi5Gx
kOw+pp9Y7NJkm7HbdRnGSoG/e4tQT6QRbyP0zdVVqC7mRN1E4YsvJDoN6RZdMYhC8mJpsNo1qkd2
ep+Sw7JWcKnscu1fLGGCElp86DH08J1waVHScu4VQBa89itdFoMSbkgEgld6dfdxJijxr45Ls+ax
omJmrTSBMF6vxidqzO8hiya6xiIFhK0p5LP0UodC/GT55Q9J556NwNo7UjH5NGRlGO3qlMOrhz+Z
InP6iCiTmfHrQiEmbDPfp/TqeviTlsRS9YUJhdvJTH/ucuAlwuiwqtAykZys6L8EO0NeLxoPWVVG
w0frVOLyfRX/DXJYFNiJWM8ARK4yk4tnHz0TQoc7Be/L4xfzh+HjDcpz2/awV1KjcrO629b+Pv69
FZL3pTY+EA7iQGvR8yTYjNLGNVssJv3/DXAc8x0SpA/l7AgwO1AVwoWU9/7tGfWrkU4AEIrTF0sn
3cxXj0VzJP983EITkOZJV+t7U8qk/BxGT+T0Z2vr+gCIzzTVHhOFYrTcNiwox/VgY1lc5N/qNZpv
MQHNlE/HYQ+XP1fGQ6qPJMpWE17Obpmtj97iDewmSrEleD7k2t5b9hRBvzXat0LkO6eWDRMRE1Bk
eqmMachS2EjbXjlRtUU32TKT83F0Iv32knIowiYq0bqdkjwwxOf17dKQZNTnuS2xAumPJ2d7UlYV
mMvw5xWwC3hVjiPdAbl5EuVddTR7Xl82VHdPuvWPfrJEeDD5xzRb3egemusqhhkk7Qge3JHi8Ho9
ii1Hy5Y0b81TFGRLBZUQon40O1eMOJhMBk0jHV7AdhRsPWexuFQ+L62Y/Yw/9y97oHZ2w5IEWeoI
Y7VbaCmcqXsF3LyBD4o2rxHjwdPyF5toZa3SgZtUpqL5lSgIFd56KcZmWqbQpZJR8LhNhixchihr
3gtXfen4CIcS1MmcbF7YxNYQLEcJujE1yovFSskuKa6lrmddl4YhuCdou01DpYNyAexLwMSU+Wxu
5dIoSkosiKi+HyR7+HW+EQoNGIrw2L2YIFOuYVLFywEQK08cfQ5vGrlBMLvqRgotjkHtI9etGkfj
RN0cCprJu1MMIrDq2hasqpFgLcxSpw7qgyO/0hCRtDm7BSCdMcJHeqnr9TP8STJMgkDNfYbKlVE/
FUYXfMovwjISe2+62I4inQPkIUjso17Y0PCN7iLvknHL5u8Qj46lUl/NptXqxRrxInAUaI/S7Y3X
jbFaTaEyLZ16C8SuAzO5MEuO+nMJYe/sCyYjJ9kWaRjrXJxNz/hWjNLeLMmUF2Uxh8TRkFKPCSX/
cZ8ELUDSykPZoViDOS6iL6px+KeHA5gJeX0hDfEVi7TraIpNdbD7OZ8T7X3KCPLWycWpIY3il0Wo
cCRyg7NceZbiufYLxnrbJhIl2uraTVsmO+o/LpleEAwFCzi+UtnJpnVzryRBOujG1ei4rbujGk9U
aebcgrz28nteOUwudmJCplmskgSJCFGHxGPM6ffzind8XsxRAnrdXh2GOh9et7AzTG33kf/IhAiZ
HOZufP081AiRW/LlC9UXy1njK1jj3geUTJw6VDMXonAlNPnwW9l8WNRfaP8x4L8exTIhcUgZdA2v
Iv+o4OAlDoBLxt/zpQ6FkIkw4uo/4QfnEId4MtlnW2PkOzH6sPiqr9nzkMy+dr5u2/KPBh9+yzGf
Bb2QCpD1qGPLp8Y8SuVFJFdxW0puR4sLGrKarOlQDmLSnuPjNxzzLqYbPtfjidncZ525KdjkWBLC
UF10euOwKgrswqzSz8j8wbESTLZQ8MOaWHpUSSv7VWqI5PlB6yPi9VkxjC4eZgFiUBGMtn+Jk+9S
CLhAfk6xvnOxtAXtWuRlaxnouevuiOaRxe5Sz+9A9Tj5/iiYQmqMUqifMEZEQyS/txogkbGu1cTd
vs1anBmzuOgMN9ybqt3CjHUsWzy+zDdbAOOOZ5KKy8Y1KujQi0uInCSdQXT4tQuMfO7c2tzCOhX7
XACOibYwg8S5cFVORfPhcoR7mD8ZQJITyn76g792Bygndo3nDb/lpoe5Cb/Ftrqlu1mrGvWTL4ux
Y9K6EJ4mQ03cUqn8LB9YQn2mwpp8TWL3ObYUYUFjGQrEa3w+FvJU3p/EFVdsapwaHDECRtlW7IUA
HVWXikBhw931AoK0ow7H5lLEgn1826bYH/mny4hBEH3GRj06WbEUYf1bx5lZFpWRWmfTJ7oNAlUP
QwwVnBlhHYUPq635nrPtZMxf+lbJ1iYWfSTXM7Au4ZJgB2ag0+NEgStPt4qvC6Adt9X9pCyDKags
aVasyUB1OS6UB0ScTN9mW+QAGOpOYG6ixpiMdky2WDFqzDaBuGq0SDzIKkW+kR1viDY01jbeFh0A
rV8mCTzEg514pPm1NO4VWDfCOFKlIedWbxFO3fDNsxOY/39ZNDH1vx+YOjnPrlw2R/U5HBVWwHuB
PFYu+qAfjRAbZ7o4bLUjvaUXhIX75mLPQyRs3/XWoAMJANugXWOQHHyaGDm2v/M1jwsBbJBhz1a/
14RpAEqzCgnjntHBA0J5mhRM9/wKYsDe4gpHn3l7UzLtJhQv15RWVZsBp9LrR6zEfZlt6NKqgpnV
DxTAZL9XHyFEDuKcarC8fm2sD1hsuI+3M1c/1z8JupqYZc47sm/qpEeyIVgd+IiSyM9on5Eb4TgK
MUE0N1Gop5PkklMZrdYdvugKQiqyP5VE71gpUMkliJhkxCP1havkSOWHEBn/H6OfP93PgAyDB/BZ
gew2uIo34414916jcnIK5Otg4y7i7VS6lOcsUyQHI2pipc2sfEaWNh71/IVjUaw6Dx/SZRcrVBSE
rDavrU2MdKfhrzlPMuqFALAjCXCt8Lw6iCvfgAbtvccT6NZya5bEzNJFcy5halLO/I6JXKywddmQ
/VvQlSvSl92fcZGOK+jneJbzI6beVuPt9BHiDHjb+edMDLcWT3lnIWvqP/hkRx6X9TDKQvQG0z4F
BPId6HYdeEdui1tDn2BRy7PZvRKjICkwiMBxH1PFYetRNL9EX6bLZlejEmpe0RNp2V6G4xxBNq3r
xK2zT+ZGoYhWS8CS9XrzEzsFtYFEgkvRyFY4zTdYL6jw3d3wr3F/Ign0UcmRDE6Gc/2uIiuuwxaE
Lfy6yhoGBi5NiXyAPMY06HfagCgRGlfBymLpjaH+KIVBI40iYjH3PAVUtSoozogtHMERCgLOobIm
TYNxFMCgvMkZ6kW8hmdZaO62fo+UcPVEzvz8sb3DKTRxL2xsTSr3C+JlzOPp4dX7J7dlmVDyabdj
omDxbju4lwhnjxk94FF3zMIar8JDBR9fxoXkHWQrsJD7Gckqi7xj5UpaC5PoTcf1gAkPIfEERgev
J345rriWIEVpJ+gNxAY0RfPvYWyg7hZcsMWgR2vgxNHvnBQUEH+Kj/75y9eBTHj1pFcJahYAzY73
zojv1udn3VcaXLlm2OYv47Em945x6xv9L6D2bhmNtVprg4HWBJGcQdEkc9mY1lpyJzMc+jpxcGHB
UaiFStki7dL9jCZiwzJFO+tgLaqlQfqCTdBWR5GrrsmGzuYsbQLwmmvVK83tPG4QZEwAdGlyfU5E
D5l1evefgrw3D6+YwFkBcXNSqFpiGmQ9ucNdLbHYZbk5Cr6Zn94sCDy1khRDlMNnvkHfxolgDDyS
CCPDTqiG4i1lY0SQBfOaWEkb/i7pjAJ2CbDbGEtAOKBxfTn0l81JZEJ2RqPMpIKNXIODOiCg1fPU
gI63ioucu1/OjeQUQPWDKx1LibALEpbWtQ6OV6EexkKlByp2/ImtGq5rSafxXLAwSDxf9J3/pDtT
I59f1YiXEaXwvP5xssB9CM0fw5j3dv2MwaX8ilQHMqR4Bl/IVqECkHa7gEdnRGfXBjra7xG6W3Zy
LVyTmYaw+g9xUb5t126rWWT/O+/9xwAd3AZAFTCuBMCcr6j1UsIn1Gd9Kz1JeBh/mIqwKLmhl/Ot
TxYFFRE+DEA5D36yD6T/1zaAqjIC3AUMtE2DKdKyHxCtKnx2WhURnHs9BKpWFwg3kmWUsdCB37YD
cLSwER4Q+H4fHx3iD95/sPimW6Yv6KosUs0Cf5s3MDaeo2/H+vZn4LHVcPtgpCpbJVu7senPqyBR
9O76INC+VMtfvkahJXtMZC2VS4jxZ2TbSjoz5HmYADAypCCiPQYBszYXVzz8kqfcEYqdKJGJppGV
Ry5CyNeIGGJjURZK8WZoNt7Uhl+4uTCOjEX7BEM4HiH7aZZ8pWgSRNJdFhXVZgxr0iQuI5OUs/WR
1biB2WOgIBefB9203YLM8GSqRGQZeUAccXIEeRXQjI4p9y0cbfLxyTzgK3aUQ2VAxHzsBzQDj/87
qN2VyIDD9X2uHVrj6UQpGkM2orOGSPE/NXBp7LqNuVthz4D9Xkky+NwaLGPgmgske4Mk40V3oPzp
U9xXxwZCqaB2bBEat0cLxlvjeed/btAmFT3FbLDyyq8HLlS/2IOVGpzuarIlqZnlgegY/Vmu1zCe
E2fgsAHsdly3/ocXyQgQL881rrMQ4gpAe58CKZ+LKiTaSP18kIgaKepnXaSAg5hLrGfaYzMhIXGF
Y1p55OhgGGCsH5AIqv7L6C/0yuzhKna/IGis9tm5LODQh0TtQuF5MA4WSp9YoyY8apm4+2cKjw7L
Khog2phJs8V8oeyo+PzUGEn6b17NF7s9Ph+P3HEyKkOpZ+2kI9Xq6SwflBJnh8RSGx/PiSgvb83p
+7+BoY31EwhZzJoVpA9a3U7OtG+vGfMBOHyd/2/jIJvfZNP/vXrH5CgT2pVEJ1vxB2JXVC5/2swI
oafMjRLL+h5wbYQFq+GM9CEJsY5vRposlr5q5GmL0W0W5Pw+R8GFKjQjnFH5uwm+j6eKJg+jL31A
fsPvfQmfzWuT1MWhRqDREZT9Rhoy0u1J6ue4hnWkAPYFfjQOPj0ZTk5aRqgJ42uOBAH0PebCV+cY
rIWrd4tFexQc+KHqzoe2U4e4mKo2ZGAHuVAEG0RvJLOuWqAJcTPAYC6Qz5u7x57fgxfxN7FDcvm/
LRTg5o07t7p4qKvap39lOrP6bD7giCWCX+1l3S6ZB5bwAWzjafH/ZsU04lqlxFc60YxfgjHt0daF
CpdvckuWgxl8PQxfBeQMe/gwY9bnVTaOqJOgIyJLufE3aiL2TZKZ/qsckFbcGtcZ7cFDietu1Q9i
GrDGKXAkmakjsl01mQ19lbiS3KNq4zSP/o5Olakz/9g6HbdcVd6WymEobJtB/kLovPg19NluDA4G
Qc7VidekCxBAbJc0k2lhXAjqkMNfB1uF3I9rp4jacApDOR4CAaYPIe53ixlbkQQ3LgTfa7FgL1OR
TizqgKkYoEaxWySSbxrEyWe/SB7HNkdYjWjYsLLMl+J0kF9gQaTCfmQgDC2mtAHsvkNFjqcpBXe0
7U0Hg4+zBKCDaMf+nVFkuFd403ROGZLUjipHxAWfqCVEoymX+OOtrxsGu9jwjTQyVl99Nadn/IPo
u2XXLVUu3meHEzV4iUVDCwUD08JjwSVa3wBCBJDHyxpg6jWh5OGIgdsDHEKT1vgbPjtjitLLi+pI
7fjM44b3AUfl54Y8dda2lfZWAGYA9RvkZN0wdH1n4Hqa0KkI+GnmhJ6YPY3WTOCbHUGuKQ8UN7mV
ZnERdCnwwQMa8DYdaxOGzAEyQ2cAsiI6kQ31SDN8KQI1D530zloxt9brOW9jOvGHjiWQUbicWFUx
QtTvu8JNUe/1ePP1wx4v4KUSUCkUEJZ26sS9D4cJz+nbtRflFRIckR0F9S4iwFOM8z+A8Sn49HFs
daGxOz5NcPbr66lQdzumD80EYIzl6mG16h/9XlW28ayRJayYkkRTdHnL3lux42qNztHkO6D7S74m
FqVf72Spi83bZ+94/T3YhxlFGI52mWtM9GtbV3HjGpexRaaIQWi7zrYVpMglbcOeQAM0SOrZGnQY
aLy3oEV8KUdha+VCy70ExpYz6picgFNV9Y7ykhGBulMMdMRyp6WWvNkjIuHehfsDeL6i23lExs2K
zF2Zd57ZusTZCScXLTn1MYiQ4FgFSlziP0wgTY+dI3usFbal+ScW5hrLM6i2+eJvTF5U2CnXJfYD
w/b76fJd3Z5eIzwzfg1ALMyNdqEb6GiH1R30tltJpquiUT5x5dcIwaFLOdEmgRhjl6p5b1DQ3lVV
0hSB2OyiDB+F2FldctotwifkgTe2/JyYRKSfN4K1DYkJGB7KrURBYlUHU0uLlXBiJUofJ1xEcpeO
vP/b6X6h9iI5c0ZiF+6e1O8NzgDLfCiAdJXnY0bugLYj+P3h60sKEDddgSZdm8kG7i3GUxhNjZ8E
p31w4Yfcp6cq3YX8q7Vg/7iHfur5Ubvwr3DvUGx2PUCAC2gg/yUjXuVrIUesrvkRAP9ckcPODCTx
9NaiNJhTseDJpF/GMc4WZCFgyTQ5oQwd3w/Eyg5PFeLk3Zrp85pGcMGsy96+6BTk12/Omh0Nc0j9
NBdQ1MQSTiM+rPi9FZWML5vBlEgNGEebXJ9xlxHB/U5Vi/0qCArrHTxwliiofm9QB4el7aFj4/Io
EZxsgWhoR7TmNVLPnst/GRhZVTJxLCgbIg+PK9UkNeV4xWUuYnv1LsNBawkCwoN4wu2lPCCp0NUV
30Qu8SuYjKwcdjRCt+ZAKnG3Js+ZG/q3kU4WKNxI5T5K44ae7KAxm7aVTCV42E+2HEBsxm6dM+Cg
fmdHQU9YjivVxCUn/NOWg4I1qLCMt2q1c9SJ4Zcg4MrKGkvJjxanEjvY+YSmQshJMxyyFK5fE2up
VuvN0W7Nj5LeNi2/onA2iId6a2Dp3kuKjC1ku7R0DC7kUmTz8bRNCa8KIVPEH9g17S7kq8V3V6Dn
9Xz+XxM7YEWmGJrTpqZK1r8pc+7qiLkuNhUUY1FDgftCXo9O6dyR3FUOVbiclJ5IQEI/KIaTdjqn
iiPT1vNUhefdT3347GWh6S5LJ5CQblZCzOfIpez9FFiVFRq1dwSy77AqxTr9zuIN1TmFxho2D0FP
L/ZHuTEe6t2lmPU1Cd+r3dtqRXd95/h7LBcEuWMDYykJI+GPburR821BTgzEQT0w9FAJaG66+ZHs
eM0RqYn6cD4/EgVt0TJW1nJSRVOyQh8lbA2gdNw3dOo0BVaBPwaZ/t2NIw0QHRNCH1x4ratugpTN
EduJu/CuRVXjgIvcXpv5+HMnL1Jbw1WKleK2qHBe7sO9TNW6lQpma8vvl8bNEl2JFF9nx/4+Sq+n
uIXY/0lxrJIg6C1LNkRWA0AYU2RfnQZnHd+PuTjaFttl1XBw+qhOg7Juo5DrEEKrJMH6CfCi8GLg
bzz+g2YBJ/HzzSKRD9AuAk+lprDLOcnD4NR+3X3ID+NdEdbiO6zZfIhg7/ZBNLVtOQoOWlm6/tw0
CHBPFjDBkJNfO3vyg/cBCEn2owGAgCpQZMYmrw1ENL7kB42pNvx5r3J1zrNRlacOw4MGpyujJygx
CKR9EBRJpH2OifE1m0gVGFCiEevGqmF9zD9STXTSwfbdTMLgqIP2QN2LTuiogGdfvfzO+28wPY+g
KTAecE8T07eRopguetqrDi3oZfSEcElvDnSe8+G0BA7UbDbT5yQ4jF2xaq8C2oYBuqFNqAvDv9L7
zzbfv5/Ht7FEPbKrdopid6uqPKYzwDCM01Z3UIyxY/olkryBZfUBumR5jtVadiddX79DYSXLAnEg
tLrBkQsIaHSOmrvIH0BigE8ve5jlwmugepAgqbjvPvx+xv/zLiihLeF2oYsAngNx3v5wIfGAEouW
MUq4e6+wAAVCLAHU4ccX2DWlzUbQGP/MJjx5Suj6AEPQidnnxVnYOUInrvK1Vrh7lL6mQASJT+rp
gERQyz0KSaOjVbFnOvNWXJuybey4PIiYXQSutBu7MdKRv6aizLixOxnG3b2JrvLFhSne3KprXHf/
wuCLSAz+JHIspKXals8oMt9Dgt2RTb8u/X/GflbffaSEqBpP0I9cbW4TmzWk8iRngqIiVtd9tTNJ
OYa2McHX+zlpv/TF3H5+ZI2jZOpgv2qYmBnoTofAD4jmW/fRaOHbRQ8P2y99kg9NAo61bHAjJtM1
vV/WVEAuaWS19Ah9jn/Hoz23UmIJJQuU2BFEeDYPZ9mugRDRf7qOCB4uB30+i8du5v/oO5znVmRH
/pXIJdn+Ny8XYwv81KpqQRq7G0KsmjQYqMgNnn+b8hirzDy4Uhf7Ujlq55uikm9LjW9u+wl1zwuB
4Zg5RZAxLiLxNCvKWgEYkZRAIw5VxUx9U/ohTjP6SjVMJRY/8rNQeU+NDqZPt6ftYddVncfwr3RX
hWeRgrZs/AwnVXstpG8yj+XgCEVf8BFA+3R4avqgNT8f33q570cs394dpESsVC1yTdIkomcczhtu
UfJtW+jGKNgdi5383qLvNvzvkccOiKlyiid4315/RJq1neWZ6NLnZF7un1ItPcNQEVnJ7zZDkSCP
MqwesiHsldqYSec2+JmFI0N/t/X2wUKP8Mr8i9PGsT9vtlSbUFjxCe5N1fSkBPpaofQZPHTG9zeV
7gJ1czWH7ZMZOPEPf6c34ECvbZhom40e+sg+Yu1YwDmGVoIVHGcUVCqOC2B1zgbBlVO6wuIph8CD
V/xs3JXng+8PTEArEhKgWJXwXNZICLFSi86Pn41jlB4bHwIcTX1uDbJEpMjqZT8I9WzLPOfwbsEB
zZ3lndxLot13R2bLLb5SCrNi4QXskxecNHHupIvCnSRhocqPyVHN6GylIav72fz9Xsd5TCG2lGD0
Fj10RfbMEWoypk1Da6/enUMV9Lo8BYkDmM03W42SS0sdMwSRYHag+Y+BBGacrEKPlHrFnYxE0euW
zsmW+2rx48K0YyYTAQKsGaCJumzH7qJDMWOxzL4Y8PvMuLYRY5at+bROZrjAYhrBBA0X4kfZKmxT
sEEKwDUx/I08dULXTR5IFFBRRLfdelMxi3VeFCG2n3IMcIGWeXJiFv0fWhDTlqOIsas7/vAzfgQZ
Sh4cx1KKXDNsAm8bRrt5hPaODbDlGnk+hc2ba+SFEuovy1cgHX4ciLWgCPLlcRI6U87i2pTv5jya
dpnnX8ZHw4pUPeqrnujSPsU5Xv7M9MU0w2XiGyEWnJLqhVb334VaXwayySMIz+RtyOwPL/17S3UE
hoOl11wimpIzf+Y4akxUqgsO8YxUw3+tp9/LujcKZ6o55UYisapdzt673kkUEjyxzmmJgnmZ1f6U
T/hIKSee1I1BZg/cLMYWV8hvHvpyv7y66TwaPt9Kw64jIBnrB97E0hPhY7MHk10S/LTyaAEQUwhx
nm+7YFRRaRoe2oIgoLZ5wLW4Djat/f8lE/B2Vs57pcEHjhA89spn2rLsknHh/WRADDpn4aS15bW/
2x7o81DTk6jL5RGtq3x6+bhWEvJ9GmK/VXFaTi9bN2NWGcEs6YY5JtO5vKEglUYKsHPhq+Ewqo9F
Om7F7YusS0JHhimbXaU5oQ9B36E35Tnok9Xzj/dqRD209nVQq+hriDKHF9mTsTlrljfhZb41toBu
vPOAbBXxGMwS7mGtJ54Em+o6UnovKqSgF/HtLd8dytJ+sZI3761CLSQhF5i37Hx/GSJMq/1L3xya
Kg0rr1+EIFoJqVLDbmxX5xC8OMy4xTi5uFmFDV7nBO16GSo6gbqMDXGYIGhwIfSxriyycTtOyXPN
k0VzOw3PvGJRjOHyaqSyo6KxB7Kkp/qb2fx1pwOcam+qb+MIURB/pNpf4pP/5grY+rtJvHQK/GLG
Ag9ivbl5KR4hexTxXKA27w2i9IyraUtmczuvOeD2nJ6cwdgwm2duEEYfePwyEOB1TUiwcOg6ECer
QFWu7MioGQLh3+wb8jFStZVoNlQgbKFyxcOlGVuWU+sg/4a+atRxPKWIojHLYn9aH1qblAyzrAod
9x6eNErtKMBVWPkr8vo6MI/u+Nw/zjXPLdrSBrcJxcWf5rlmpnFgRl+/P1/AL9/dRlrpmqYHZHq2
7i1rAHW3Py75btGVd60h96dzx9CQeteUWc/Dmh1DMvHkSKd4+ghe/C9x2/uzwILs9JgMZE4bJy/L
5wJwAe+EL97baK4FqxrGOBfhuDOdqxWd2qZTvY5qLIsW7Qi6vGjqwo3LLykSbkDpZiTYGgzCVBom
W9owzBidJpE2ykBl5nZhn0Gt+gqzf8l2lgwyqaQozff9xc6Yjv8XnXUPrd9f/1GFYfbIZp4L1kMf
BDCQhk7yCd3Vl5qovV2Un4HzhTjqEx+GTd2h+1fvftt3qnQcZ3QoQaP7d0nk5tLltHTP/Z/WzW1G
z6ltVXNjXI5TB9y/8NyHuBDVvzwbOv/n6VlltgmdGKG9dyqwxoNtciK4y8Tt6Ddytjm8yx9slwkL
FNGuXAkPPQ2/WjCCxcEcJalFsxKNJyCKMAwTtQNrsd58Aq/JycKNv0ymvIaU40f3Yuu775gJLn5V
dySDQXO+KVskYX9XuEm+t9ouKjXklcIea7cTZL5wHtMYKs4EY3Q3oxaUiw8AIG8SRTCsRd24Gju6
hk3PHSGaDEpto9rvVMAqRJEjgiArunIDjdiv9tlDyqjK/i1wRiWBNhuxVJ1FW6IWFDSpKuw4zRUI
BIBNKpQrBnRrECAab+8N84F0I3dLjhYKt70uN+qhTAXc8vw2xex//zkHgVu1OaP9XRnhZYhLP+nW
NaLO2OoJ2vzJOJtP1sHwQz5RR1wwoUZC/3Nmo403mOHt0FPZXZqU9UMyreITqPoZcBlvjeEcItH9
OMognJGeAminrPBJRdr0pP0eVq81JEfwJ+Ib1rxNPSsBbqJ/H+ZZAbmDUgw4YmfxM3yDQ1n85e/S
4/jIGNLe66G6sJf0AnRTJz3dNrzWmgyt6BQ+x2ue741sstBKdfoBd1F3R3mkomR1ciTe/Pc/p0/j
wiyAj1YtN0MlenjVzimTccX6/IsVzfBOLYpRAJ4cL/5D+2qkEWAj5nzIpLhNYp4xEQGpdRZ4gyAQ
t3lHUnZACaAm17raf03qqIRT83cmMo3C8CM4UPIqZOMbUdi9RB6JT/KDLX3OhgoiGSPlQad9eAxm
5xKDkDsYSfgFRZuzoubfBu0J1+ZxcXK9wKmd2q6ZDqxCmuMKHjb/49cSSkpBP4USSf728vb5kq05
6j2spyW96GHHPlxaQXymqsxHdqd5n999NmSzPY2+FK8hCP4TXKlhaolWMpO+wxedlsbn6J4iLzs9
iIUn7gSo7iHoiTHzeI2mS1mN8D0vOQ6pkKS+Bb4rYXqV/NugfX/lAOc0nk4gFLqqxlULxdgO7+R0
1kA+gS2hjQRHAByqs8SWf1axW+awK9XGp5ASWYMRvNTt6w7YXRD0UuyFy8yXdLwxYNPLkb1HUBn6
jN4f21ZSaFR7hIJgGcrfKRRoMbc20tYfYOnXEkA8mjHmSES9u8J2IkHSycBZmoaxeW8Cq4GQiM+M
kRkOF0NpvUoDQCf/e3HzljBPCNjNPwVwTbFNhPamIjcRBr6gVp9OAl+i1dO5OeQh1tm+HoRserbi
dA+u4f4I+2wadI5simb4/SaLNhUnG4DFq5ru8fTfUU/Y3LTIyTrDxsvCZ32ayLBKPIrLac7kmY8L
iNSRpSLh9j6wZwOchE+3S+/Y3yPRnPPvoG1JlFsS/Li1qap57VWPf2Th/wBRE+uMmH+6XeWuJnMd
bUsrU6gDcgqRMhVnwhSQEZ6euov+ppfnugjQXW8npIQWu7UXyrgVPB2mPT7a5TTP6bkzopK+beEW
WycfHUTQrJmk82s6xpALXdLddZsgo2zZ2YW+m6HF2QgPAHa50hwRaXKArWZVDoOYthxp2fiijnPw
yFmQA0pDF3b1cBjKCgJ+Zv2E8HH4R0/iv12PFv5JaG0wumxQJrVMJALYRB05ifjBFg2wVU8g3um8
KznDFLQnKdxhZOmx5UFiTbuEf2LjF6CVc7ArQUwf4mX7XlDUD/vJ0/Q2Nn5+18Gg28o9eZNmpG4u
0QHy6oBoTgrhjP1bzDePS2l6Tk8zQXQ6oTutm852NjBbncxG+AMfN1ZuLAdnflKg+io/QZkiWtWU
9fBMonQGvQpiF7ppqBydrIoI/2MvnpNlSGu616WKfa60PJqV6MM01amWH0afs164eLWiPITK03I5
2QtixCmexQzaH1aMPPJnqz8IZsZE7oPf7gQNNEZj6ow5cXMbUyBcoGatA7DWXPIN8KaVljTFY1Rt
56wRCWnKhZ3DvDqGHD1dh/NaV5rydjgak40s3t6kKgNLw1uycajrJXs6P9condwjXsQNMI5qZ1Kf
VMIREtIV4QQXN5W4dMuioQAyJ/c1A9FCk9Rp5QILw86QLXJYvRkV90vs3mS1TJ4ps4YKOE3la2d2
3iZ4565n17RM2d0AZnWdgj7o++fFa52fe9tQcxbJqAlgFN5gBFvujbHtp1LB5Z+E4O/lGZ+TxEr6
Cpk5FCLqeZzc+R4vheIqa4x98FMluekHVLRd6aoDIWzZihEAyv1zpjTfeR9K6JS5A29/i7KUz/BE
2xddckssN9GhNjjeEmgXcVUYx3zAVUBSzec1tTod8F32kz5oYR5eUHDVFKVLrMHzWdCDSbC9Se05
6RFnOkAcgWfWOi2hR5nKKohu91nR5yKLFvs+81L4m2jDuweM5PLR1kTxle93Pwy3K94+aBeEwKam
rXrumxA6ZMfH5b88R/7x1A7s6XWmq9sS0XZdBqBrNLEBiyDQ7PMS3rdFyxJp3SOk0AhRuUZDq7Vy
QCJ4zxHfEf0pXX6gGO6vPthcqFjx39Ti3UYcEFofHZu/h0dJP3EaHkkzQAmViRR2BJwEuHB0wLvW
RlgKmV8BVdDMsPirC1ZXA1wrFv0ZVGtcopsUqKH4ce2jVdKyNgRZiFWmor4e2Ai+D+9Kllnbeea5
cOJSwFzx5DkbPtKTtLctBaZV5XmxIaJIlEAyWma9uUT6ixadlyNKIEibCKy12qyd3calOK2wO7+O
FJ6UgkSM/7eG7dXpRmln5s69Jt3jPR9mbbVdciQmO4iNOjOVQ7AXXEGfSOzSrpo3JIpif3MnWdEs
vMsTV52TVUsI6Xb2bEKKY1m71FZ+jE3PX1/rkNDJz6hASYSBDGDU4AC4IaXeLfwcbBj4A2b5BJQi
VKho9JDzCCgfB6gupTw2c9IlYLvlUAjommuVYWKKOmLCqJSDCQbYRYtJAWx6Gaz0C9FAd7NfngZF
SRQ0qlKVpKvY45BK32xhGQ9I8PDA3vPqsh4g1PtryGcyd+nGiZcwlKPJdLgtky7rvD5MwlS57Uzr
wSmWvlVlmkbQL2VtLJp0F9E4zxgYiYj4q9n6i/K1Fn7BbxwFwAWPXrWDw6fvD541m7tNS85YinOg
UVYsskZT8zrKzlfGjQtfDD8fMrHZNaj8s9g0rLI3LfrCm4V8Ye8X+kpJ9u4aiUy/1M67Z6OY6IYd
Nw49HOX1xLoqZj0crh8f9LRbJPxAEapoxUPzypPca8bMrmnqgHn2zS7byrWHJ8AKX6uRa++/f8V7
d0hNKDjCxVUvtLohwHAOArfNcOtG/EvtoY1eKhipKS6o7jKjBqxCcv9xNcrzUBJZwfNXr49bibII
B7x8hc6KM94t/bSqyWxZGTU1rQKhWbUn7+fcGYy/KXKrvGRCTqtjW0Nnxbuy1J6m/2iUDYT6SyYX
ULvU7UOj7/N2TkrJ/iov5FWwLiFEVIW8m7HBaBddCfN28jQClxqvRfgloz45CyWVIDqBL//11LK0
yJvJHwDXCqw7brqlg+pKMEfbV6WyHAy1vMcxZ+5FyxKmh501MZB5aQLqDcd1biC9c5CRlOqByWgy
quFcWHbK83UmxAXbAFeynOZxCCg4eqZm2GtZz3s0/DFbNHUIOfrFRQyN9mM9p6qt+DOYAg/O9DPi
bNGIxb3/NiF+6KNOn/4spdQfvdt0+EKVgs/i/3ynVoIm/jKMWmLXiQ0ksddIUpdAcf9k6vKg7a9T
UftcNe6EiM2IvUQTeDxaA+lntgz9eQTmpA0ElmBvhtsbvOquo49El/pwYf93V75YerSq3EON8hdp
ePw3XAJv6MppfZWJbKr8MsQNCO4+YWbxlUCicH38tSP9gI7d0Q9w+tvo+UU/q3o6w9eKgdPVF3kd
uVHD83y53YBSsBol2HaOTYwSk6cXdZh5s2cjPSJMnJxfZD9JAOsj8pKJDhnL5S9B6l/Z0jq0jcZA
ijRuADxj0bah8KJ5c106Z9+N8q9Gex+1+Wggfbouyg1XUxc+r1ctV2+K9omwhT+OXbUZm2r+D288
wm43Xg+LkrxncEdpB7OK+lrV1HO4IKNNL75FUfLuVOwgY8rTQMSIMhJ7P5UOB60QBpDNHPHLjaEF
bXnoh9w3jdVVsKmTSR2DNHsnLcvwBJQhswGsgogC54NTn0Kqh6lECYCgBreGcikbVWixmlzhZAd3
+0drvTo7rYa2jNEjSHuViE4q28LwtUaCthii+BmEicHWsg4URPXS7GYksvkXnyshsQJdgxxyW6C1
0WpmjL6JbrkFkvQ/wl7aJ+rPBDR1VQnHG9f5s/MR0OvpqSIlo/JPEhnPkAnfSxGrnxTBQOS8GEXb
0f+f/x8gQcP7kt6tEvCGt1BzuGFffxBCkagrAVRnNCa4mXEp1cVfq0xVme4sot9m61lKt31pY+qz
VsdFf5Ne7mpPMhzmFr18Zd6teEDwMCJcL3dsVGBm/0mxv762QbZJaKy8vjpnbiW99W+6vmmxkKXh
ORh0EnIRuh6xC74ZaQrhkPenrqAy9npEJASQ0FIhL8aErA/Q5SrvNU1Xl5sSSSoH8obYdYocP7pG
x019GaUS3CyVhrOGrg5dxpZYJRNZIt5eja8D1I+ZBZiIrnRTfVxi2Ii8kWeH6J8NMj2tJARFOKEi
4eR7lNM/YQHyORQu0Kt91f10woK7HHmvI2h+ff15sBTa20UxjhdqMfbFc9mtsOA2VxAICOniWRtN
NaL3jfwNQVaMCJNLmoHIwZBYrKBEJzonDiKuL+0F97dVjsmJ4bWo0pwwqQc3pu4OSBRnkXjf0Gz1
QWmD/dFZiMf+PGqLE4YC/1ABtX61Joh2k7WQl+1z4Ez8VPNEhCJvygfLYzub4AWK2nPqmG5bH485
5ukZUSayp7FZJt5Zj3/bMU1atMHYjjvMQgVneGouerwuI0D4fMoepBqWNbv+nNB9LMagEC7SlG11
GaIKhIGjNCRj+fQrdaFfmDDL//6WHJs2fYC/RtxgizXQJ2uFcizuSpHVOsW7O2jCdB9HztSyk6+i
LugTdBBEaDOnl2cj+xU7lLGrbDW93w05CKQLWcA+XdgqJ3PM3mIr4FdwG7Cku+fxB436ayhwbcDV
8cvI95wufhe6m6pE0nm7hw8uV0PPZHUzSC9K+PcfIxZ67idnvGObVoYYR850HE1jl15Iz02DvSBl
xiCETKA9WrxdGlJTd2hUAI7BbXA6zZAOc8lbi94gB9S5/beB88QNrw4ET732K5Lh8E499EPaoQ0D
SR4VjJm2EyBSlkCdfQS5TNoR/LZedv6wZoJjymxcQczNOsamicJeKYx9plPqX/r5zSARJoGvXKJF
Lo1731RaXCvFLDBx48h+UTpd5xr9zp1u/q0tNWfAvx5b3RBqW4Y16/pV8heYbwMc9UkN+YOvsCEt
JIeNWZXWUWMz5uscFewO0pNpoPc1pWJ2gbU2guPUg5Kd9wczl4dsDDKpPK2WgLODlyW8tFgkEUm7
e5LUBd3taIWmBgqU/RFnND7kCGzSnab5JHEdoNd7dMZRpFIgoOxh1l57t5vsEtjf0vautnwPgL+g
FZL17UuO8K1rfOl6j3+J3Xim2t5kdlNltBCA5QD8URDejz/TxQ5QfXylByuKEZwSIjgi6yjpdbfi
bi7hEIIs2c6Nc8WVUlNfYp8X74cbOvWKG342U2twKvy8PEzulNP7h3kG+hAK3JcP5i10Ecl+nEl+
vVIuBYVeHEHuAaSbiOwZYZzk9bO3W9qdGxxr6pZUka7ebeKJDlfv7no3u8ijaDue38EKUhbAf6Bm
dklhGEg1ps6Q2S55kWQXI/XW6tWmf/TKXcnjAOo/vlcmnZ7o3Hb4rvuT7/O7d7tSI0HnCBl2q5I1
hRX/mwCLWorNLM45fzD3Sv9ACdnh2ZeEuJM772k4LxMzRZSdI9wHeBdMr8wn9MOl0bgsCpSiY5PO
p6yhiczbZqDrglnp5f7y/DgxSAA1aP1rHEAcjvqbuiQJL5ZaSQKBfhyjrVeJGXu3ubNtMjO0kaJ3
RVZAa/oXwfSu8GR/IaThVs4L5SnHmeYc30SQuxFPZROeBQI489jB/6LMpGIVKjm9Li3co+TTbW7j
7CaLSX73ZqJrh0/L3UKJh3xH4RBH3raIzLhEQ+mcmhCajYq/kChJjXcl6iuE1O5Trc0yZWaQGP+c
82lRgEaN3L5gGyxQktbDSqUyNivJHYmVjROqf8KARzhBfI9Q5VZ3KgzvY3/kB/rC/9gv1FJRjfvg
lDB8EgDQ5dLuql7VjceQPBLJWG+udlivEzyaIuqQW7vx/0dOkyvCJi2ytp510Z1nJXtvylw8MSbj
Kvx9nGU3Ie/cnA4Ln/mLau19VgsWy3PtPk/C+RN8czsS342RtRYIVGq+YKR5LkFEEpF69D+Mln1O
h5R8Q7tJI5jHIz8/rb3krWo2PC+ANsvFhgt4Y3bq5g/CrFIpt5MxCcnUQ1v4DVH45D9RGqwfO6hu
W6WhvTp9GEhFNitSEgEExDuXZjCEUFy7R9v+CBLRILj9dvq0GXkakgLhCPooUiTG00jOjAiKfRLq
6K3u3Wp6Ria82np0VXdp3wvGTHfklfDvIsm19Uy/kaObObr8bRhEqxHa+j0jeopOzKt+1fWzqCva
/Uv597Ox6Kfz/NnTwr5IlwxyaXqHGpYzdDZy/l3syYfp5Pa3+48ZM37EtHKBgMneTz9pa6HswiVV
oU4LDe7QXHdMRtnnu9utuFB3SpctTqdtcXz7jCQd0EXEYWoU+I17KHGV5t2UALdPXE2cQ/SqUvFN
eqQ617klcfh8kXzx1nkrzgs9uu8mSxctQ4D7Xlb5q20OY7fu7j4uhXo7p2xfXgvrWHlOJFM+r29S
l4tG08rLZVqJWMPA6LDXc+86u2bP0v3ahe1OvWeUdEBafyuSWHHmPwkbF7IcqKo/mg4RYjFXKYSo
fbp3zZBnYHNuJhvqcyoiTbwcGwaPcOcRuXG/+hKDOxOuJkwk9gFnZvTVMyFriks2DoU9sZW2xdD8
KPidxATdB2oh02jxMshePfsFJuJj3jkv9R42tXSYIX4QEV7+mRWD2woBzhlxQ+F2w20CDf5NB6ss
L0i8cLtWG4DCJXRWvB/+pI02yYtBWZmLpONvdY0WIPMdf+SmZNiC9TEAaCBkrLm/QJeZHJXp5QII
ljOtxbDsHAcgE84KLxO1pXLSgWURLraKn8z87PyI8Mx+sKW+mswLF61U5tnWkmrYXnlUmKEl7MpK
0tcdiR33fTEjbzeUR/bR8u6VFSnS2ZZLQ4cUsiIUlf/wgSLjnbKk5Uz2auVjw1/2XziFA9Kgtgh3
0nqWS2a8o/h6vc88ib6SxEhIdWLsb38Z7/ixS5cmS4c0ialM9uAcxFNxEC/HPLjsaZWK7bXr9Snr
EDa2KUgH4lhpV7dPlAB4DY93KbyKvzEXe1uB0yJSPIJrlaT33Nm89Q+AA+AvW680T7s21g+32NCh
6f24OOT6PpyqtuAVey8I27GzaEn2JTlYyzeMtWz/IPMM6aLhzcCMAz5aqSk+JGM6ssbmxG4/QDQI
wg9YDDejlrAWw2Z4f8exJN9nekzfecxp24nXlyjFjhrujIzxnikE8r7EYTIGjU2lKalegHLFRXKJ
GF3XtS4wRJwn+s4Kg8CxV5m5aFdG2Gm111QaxlyoFieCY03D5qkg1lOrFXZ57ojNKLkUBeL18lgv
mg2dtTupnx7E2rYHigcZI1b/tPf3UUJWaQcMTOYFkqTLxMBWJ+LPZmTQCmvuoNIJ+fFFM8uRm0hD
0XbKudICWkBFlLxlB7aA0Xe2pKFq575RwJuDiFIuWBqaqoCYBGaD7Dc1U6MjZHIZjC8WwP44b7OJ
wqW87Szg3t8z2c2MqnOwDszXN9+IR0yzF5MxeKDi1zvBqRUkXZbwEnmKpCMJ9x09jaxq6Cy1UPq0
cKHjaQny3POVskDQmHT1syPES2yl7H6rROPIcUx37QujPk6hSYkzPwFzaAdeT2iFlP0VfA0x4N4/
9pJSmJpsmHpqUl++TH98d4142nRopXc14z2Cl+w9SEPg1QovbOVBQwFxiCx+s+Z1IZ+tl/hN3v88
6gTuevXMYN932Fqh51hCOeBM9XKFWsNXNzTY95EZUHpazDYuJ2RnK18fMLnUydVycsZ1PU6iVPXn
diI3+VCIIkV/eu7TES75dA5kTiPDYt5liAbvj7oTsyNXKHHozslogjV4mwr6AC/csnZ2jXueFd44
SzSa+6uif9SiE6TzBSzlPu2cK63bwbutOhMV+XH7UPKXN2ogOon/Zj9VK06xr2Nb0o5E3UrLvuci
EAYJq2fuhX7il5cFJUDWiOujGUCmTZ0lH5ZBhYA9w6aDABfB7MwAbVd3EC9vKKcNbB5k0oAG9+NF
NVxwLphR8AleryIzeZbcOVZw7R5VfHDgSm3xarry1Mm6KxREDLKt5FjLAblbS3Ja059FAcNFce00
N2iZIDUq2dIsdavE8k1ppArBR+Rk+tlqkV069VxmYw7IlYVgrwBR/5EJpQCs618E5VRi3VaP9wDJ
3cUsjlP1kzCqOGLd/Ixa9ar2fdsnhDCENMVMBVP/lUzgkrK1FopPMkF6QXZ9lCmANE6tiEK5nr4M
Lj9s0TP5gj7rVr8/QHr2Sxg7dN3lvSqT41Ptn6I/zsyyJ+TEYuxtD8hYldn+PxY5OyBvvdD6AzrY
7QY36dGSBQ/DME4d3hdOMedzqf7uNqduYw+K2Yb59+Juv4jEDpfUbquZ494LyjoOjy6kK3MZ+1YQ
T3llyFeU2G1CF1/ch63Qla8kn4DLhczVLn2viTxCuBYz8/HoyOE9sVGvrtlrkG40qmed69mlL/HC
ZIuw+bTp94GPUCH4nRAnzBviBPq1E8FNyqlGyUkSIVK0BJcmhIMgClDasmAobHno7yn272S6fcwF
QbEUuC6PvH5N22joij1tz+xkrnUlnmJjk+53CATQjIgUiSiiO6kRNqtVouNNIanvvGH47bnApJmb
LbgyqeIHsvm3JpB1/mn6QmeMHQoIexRzpSMZTkofu13trVJn0vu7SDXHj1IXjNcq1M18REbEjjaK
eyQBlx8L7MPRQqYHCWgIbfaiFGmptQdO8uxbZtjs6SV8i1Ax6fM8LC9kI9b7nvrhOL1tgSTTvMYO
SQGF9sGW0g5K2ViIZywrZ/FxaXgvgll0SxRGa5gmBMhsEwALkOm2tuy1Ii7zsntQ2AKBi+GoOTWq
nCiioLEbzeTPYbHck00pNlADTwTzL1ZTgbXuJ62piT8itLMoQEP1ArMVDo8G8cL8MorO5YSFs3KB
udDN42Qrw52I1UYjMmInVSeh7kINxoTufDVQB818Q64R0js7Tat0UFPhHNjPwLn+M5/ArYx87TtM
oMRD6+D4TWPQ7wNbwDH3hAbSkxIiTS3EfiZlw+UZo/fWO3yaXqnGazIGMJsX++zcVlGTdR+PvgEb
WyhtReEZ9LJxMbGxhL87IeDPKFiU+btn9M+pPhQqL6j0WYKYer5mD0tTGjxS6RY3P7KxLAP9LIGp
RrOkUyIDNz4T/0wxEGlAnLfp2b7RBjiDKTTWGcLMuL+aEASLy0+k+0yRbuZHKPAYB6p1+eF7sR8S
1YVZbOvFiGoYfnNxLZKA2Gh4wSLjGksZbQsRLx1ZTOdA9tZUT99Pc2WGDRseSpYQbNAtQq8mSnqh
XT7DK7LQSVdzk4lxbatHwe/m/9OiXUgLeTPiu4He6zGKqP/viYdEJYNANjHero+dOct84UT1JT9b
X2FAhyNHSVsg+S2ERXMzpN80rh/ZIhLFTGiXq7JyaZ0W105oxPsoXr2vv3Pm3roQ7gCMaeYLwJsz
IEKKTvqUnfR6KTcdEZbbLA20fCUE2ShopZpGBCkIxZdrzHAo754FSYmgbY+vMo+U2FcTH7pQFUj9
K6dK8+EU2/cZmSb4UmeInVi/v5Ee9Dn1ufBWlYacTrtA1uKA5Y2D5/kP+Oj5kzhvKSo/cvzDtzFo
G+NyncToQy6S6FFwfMl1Z1kNKquUpv4NaquFCwXku3WGHZ2Iw6nKKwigyex2mjDeOr26Taq9T9jY
BQL5Awnjj9lMe/ef23E3ToO6shH5Z25P5TguUY67mQoEyqjbOwbe7ECkMGS5FmuXWmZkf9pkY0U3
xmSb9+g6RxTx3uKAEIXzJmf9YiaOc1X+OhV/u0U8FGS85nGBlmKOuPSMec05GjeRKG0LvGdObgGL
h36tkvOSe/XyaKu2KLp6x5rHOXJCLFRkZ8P4LA8I6OYC2vQhx0/k4yX7ozm+NKl1M4tlLeQ5eNFf
CqtWOrmYTRGJL3xFk4Fl9I5xOheVE8ofNipcCyUDD0jx4NV2uR/BccpMkBMgLPW0JvBL4lZ+VGHm
sEolUPGpnh901n4BlKR/dj0hB2Gx2C9uNaRMx+biP50uJn2GqYzd7p+iEw7KpzLw9kUOan6w/0v1
ur7mrLQRzs+wu2tHyC9/zkDXJ7LbwSQdyCUf/Kj+41m2gDXNoiKrvHW+GvdXkWsPsjDB2Sdb0NPe
t4zIZYHNIzPeLFZ5W8TzBxI/wT2RlkmMkZEANJWDR6pL2wyBUhtAwLwhtuUc0IJ7ALgLc0i3AqUg
B1K/+yofkwjzpEe8mHZ1TnwMxp1/4pLFIWykip8zkVnMOaow4qMORFf+7KxsHLTHjIkiWFpTh9+Z
jFWl094wVzABdW9Yj5BxQhmM/TLMC/moCGA2dyUjqgaDH7owZnI4EOMasv8k+CUsYgbaNs30yLlZ
wVSHGEP4B8anPWi+H/ux83JaXaqWnToUXumafnp0mmsQMrddkEgTJPeuOsIQGAAFPmj68M9rUHZt
14uTNEykyAbMAVAXBCgnmFySL6B74opQ4t4/ZQn+ph2xKzT4O92K9bJ3xTKtIkYe/sLH9L9Qm0mH
nb88liYT7uyVgTWz4TID0Zd5PwPG+zuyPFRrcT+SILxAfeejQxnKP5dPDLjNBvwOilN8vh04EgKN
fWo8tCJADfkod0mvomvWdk1TqV/TOopywfE1Kn+yum6HpfszKfwOrUH2vp/O4jrY1wXL4xmgV3jI
dSk/5Qwuv/QM2srrleJ24tcLkewFvoyxR49loZlVLOMiYq+YRux5uvSYdWwZZxJCTnJg0cqBjj/B
vVUWXY+9zpPLjuXZ44h9iCPPD3tosc8YOPNJuAE7NxRPC1ntJffpdidrX4L+n5GezvItRaC8qQ3i
MNzrjfyMWkljj/KU/4XcW1stq5mporAb7asjHgqpp+Mjtf5X0cMUvtTLIcKoM47ZS4N7t2Ado/ih
RM3+TM9ay9npD5Yzw7N+jYsZIr925S+SpltcOtKGz5+A49P5VWA+Ezaee76YQJwHBm54i1VbfH8S
sw1cLS0xG79D7w3hBE2Rg9Em2Ju3IkScmjMTVn7c6/A8y+AS5B8mqDWAEHEp/GTfx357bmIi6+01
pkKjItL01vXRt1u/9bK/5rjAW0BwatGeF+kynewTvw45EUbZjQX8Jwyi7MN0WR5cn5ZEIU9pvcmr
asPHqVQzS7NHVGluESTR7XNcnywEJeUtjwlxcRlvdXJ98rA0OOBUxwnzrZ5rB/j6g2R9GrCwU7IY
EIEBLxuU341I7YV0TR2l1pubNbGB92srEKvSEaCcGUWi0c/iBh1DgftnII0UxQRwbBQlo+yEKhC/
xWzJa5pxxOWDRZR85h2LMz1R/gOc2po/sRgBxrLrpIzwL5xxMAlhA5vTcjksm8oADfqDgdtCOrS+
X8W6VtFGT0ryN9ta/B7m8IY4XyyXaOwnyL53MU5LlIkABPlaiI27nHLKjSPfPHwzUUKXmjCQmNLV
SDmswWoLzmdhmd557arfWEvsbcskjwlcsijUx011UOs/8uO8d1EyJqEmLjE3QzpWoWwZwEesC+1a
OG/rKJneeCFA0rpGjcCd7ZpITt3sj7MMhLNRbR+/zm1iNnlwwOx+vycxcoAWmvPJyZ1ie/2LPPB5
7kIyO8x1RgVKLeMYb1yl7m1YMx/Yaj36Eo3eaYJsSVma8D3r8wwBJiZNiPGak5bGVUcT5YFZCXOW
3sJnUVXhqPZkrkkNJteT6Imgt316MAI2sxgUOBVw+R5QIls/kEF3z60hzVJQcsS4vyB9cFdkiD1s
KeN6TMrRhePaGjah0rczrGPlHNoKqEUwoiegdbp27k1LgERkNaVHBgDN1EvcxJnERgiXA1OfM7uy
3QWcfi9ML5+3HYT7lOnb2P/vNvfhvFSaan48C5Di5uCIuE1+dz3CQG/SFzRVHPdYVXOtn7esDPu9
2Z81nyyRHYGsk9o8hMmNA3wxWrQRysLRhMuI7kTEkY8PfnyvdLsLJzjBqKm3JNPieGtqMEBMKfRe
x+Ly4K3oMfbOKVydHZNWL+u8IaUHn9D18SeS0WDz5AzTBZQoIaOxN6tvvKEQXt0jgrbVoqHYN2Ab
ridpQ+FN4mrl+UksOLDoG1rVYoF9vtzJv4k3KPCvld4uS9ikS0fDBc/BInEYWAyeh1ocSGNtkmYl
LFTtVWWBMzVqaR8N1vr3B3lcA5CUEpCQJEewqq2zePiVpVw6aZ0U7KnSoLwtsAmShEh8G0AL+m9y
5OWiIdaB/pgwXtbENHKkLYHPwFCN7je4olH8/BF9jKDYJqbMwId/nUMWk+bof12qoZcmH+hNXsYj
w7SbdcwJAqe+pvKpRD5Lr0Jr+A2jcuUgCnKFVvbl/XXaNrNAqqUYJQe4D3BAd/WeZBd/roZJIIUE
pivokOVhL/XoIpZfxhD+NTk6a0BOxSZjSfei9zB1J0ktjGmgqUzc3NAzHbStZycMysl+zVwaPk7G
di1FDJiy5pC9s2WMk8VULG4j9SL0TS3gG0kZHdWd1Ymr3Hg4XBk9WTfi9PJzJhYaCD4Di8KmU0+q
a6Xvl7snu+FdIOWofUnqxrCSVY1YiFyMLBk5DHgxssjv/XtK8NYYBWGjo1MdiXqV+uFoLlGNSqzj
m0SWit9LCZ7btGKpc90ihn3weYUzMNYFkap++RUczZdsb9sPxlex6nTUDqIMh5Owi+mgDwWYyJHI
j0lKdXieZfiR9VqvFgjx86UIeKqCcC0pNd8gUBf1zVGeuMne2g62TmeKdGSMHXdCyE41n7e48Yvu
1RPbB1QmI2IS+YKI6HxbyHcFv6I4TXJEeog6xY4ZaIkWPsFpu3mWuuMpVpI/OFkyLFF2EAhAnC+f
yzVwiXaymm2EjQoIV31npop2OGIWxDEhMpMYexmsVAx0nPWSDbddhAXCt5d/fj/+2xfxhNm2MzDY
lgoS87QurpE+jE3h+vDOraHI/rvG3rIFH80Nbkx1FOTHT7uu/fmNLH244h9WbMW/Xb5ySUoGJ/rk
x1xgf/9UWeNcv+sQAW8G4CtF80JG54Hbg5x7PIZs6TJppHvki8Fq/CysV1UIWszhHyYtnjKPy53m
Q7mYeTacCNwEpveGnUoDeTB769XXFTbcx+mkyap288DbHXiZosT8em9tNQZjp4bF+lLNGpHYeCZT
e/bAsh8xfX/gcLUTxkIYMfehsczMjnbTrh1knW/l2/gV5NrFJ4gjBQrzy3+nkMOGfbVY6jW5AEd+
nEqqlv98NK3Jn0T27gDqXemeMPfaxXEQbPnC7EvJ3sHZLs5hW1gWG4NOsVmHFUWfT9ZbwRcERv5i
RVhpnWDjvqn63p/hMWhTofqS+zirW6HWGPjiMWqaFWT2e9KTTV6eHosT1PHnbi2QrL9eQjXy9M32
DW76xB8sgZrswLqubvJRjUvN2ynUPYwEzODZ7pRfNjOMWWKcaw8Ge8R4AIWyD5mhGbk1OMxEs9rv
HgDR7HA0dd/2SjOKgnS2T7kTE6qK5gk51+wIKErHtJNv1I+gMsNnZXCoqHynoBMoHxf4LYwyXDN9
k9tyqdkPYCzGRchq0KTshNQHgeMuZ0781+B3Tqz15NixIXhbag/UwHHDnkHHlKqiAdIg1EflfaNk
19t32C2i3l2j7wH2nJEev+o+NNJhCbHm/RaGQLLZfzEKB2n+qG2c2/uHNRHML/PAQnWcgmi04U7O
SHqiIBsKQ22VvgdYY9geVVeLKsQJM3BYx5CRQCydcmeDw6lsvuj0/c67LVnBfUPH97kaStAHGtFr
V71LQXr73H6dHvjaMjMZY/tu4Mb0VfLinZLAOKjjUuREPKnmvURUqEk72OnbfV7glqGJP6iuR+sx
5/oA0dlu7zOSs6Voi5Sqia51qHspaoeQhL35GI8CqrZJjT45xcgTK2t/bdyFsnbvsMxOT3KDQNpz
dmwWGXBVSzDYvVy+LFX1loH6KpdQkQQJCtbQ3AcESDAUlEpnhXV98rKrUT2FL+D8WYxqjBLZNByC
euhdhgTyK23OS0lN6y4zj9HUrL4jOHhfbOPIkUMY/CqzT/mlJj85XjpsaUBMI9HGaRT568Xd2yga
4n4AireOVKYK78e2LgF/ObMKPuKh0SQ8dhsmK2qjxuIbXrTxDUM+CP1oJAhPNFZPrPRfvnF4B8OI
5gllQ2c+zcgZrpSTUYg4Cngy5p5qtXjphdMOn+pzZesULc0NVwcW/wdVVEp8C/i4UO2hOqOqvxJc
xhRH5o3Yim7YC3pepmZ6+BSgBW3g24qElGzfidVKbs5sbqtP8xpJsDOennfHVkEPXKRvUHAYk+op
w8NeqYVj9wG5gBP9xruauCm8GFJUWBLYo4u7NNj0tGcq+xAB3a8vK5IBgXO9bjXuFqZrlUue+F4P
IgAHYtgsPOJQVVZ4iB9jgDMwTk1YfE+l5YMDy01YB5f1LpHCb+YjtZIGC78Zq/qi86ms5hdgZhel
icIgu2ueWBmuEea8yyiLY1vzFzKy684xl4GwgirwjTTT0vG174yDfc20cb7ULP11ZcIIq6OqJ+JA
yN7aeq9wGHCLDKh4+9lLK7mqdDJG1jzNrDex3gxG0SLbDy9d6/p41JTLrAaNNdE497KTDp18rrlW
Xnzjp10I/kUzAixktnHM8vBV1wejhVJmR6l7Lv05OepKHQfD9oIAgoOuWtDTxLvZPxlfPSSA5cYY
3hwuBR+upvRMdZdYveva0u7adrfhh9elKFL4zm2mg4h7YyzI8Khx9l3quyZDRI2R+aN6PmtqflhE
Lm+o8f6n4iy0QAzigPELTQov18DTRvJYw3/FFD0EiSUrJINgpVrNPuvhFBO41uDGRCZV90YGUarH
xEq/uLsEfaS7/xGarnvUABAB9N7+64jpGWbVoChJytlEcKtcE4bO0BKQODu5Vi9zOJGpuLZm7LwR
kG79yii/cEMIqPxZTrY7f67VuEPt8SjSpPnYxTHXra/DlyWIZVLKDE5mZcLoLeG6MzozVWWb2DV/
ikZkRnqRs7EaXfulaJuXRB1OGtU8W+84T6OJtePRy+zi/vQ0XuIlaK54p1EG6X0tLbfNv+LsNhPI
q7cu5zw9OII4RGl98rmNzkZ+JZPC9DUvkcrn0+Cw8Ibjq2Hb57sqc1TogFc5K4djj0D15a3EIyJq
RDbxkf3eb6GGKvN47b0UufvsHsummWt+jBROTwdBsZxOOaUt4fAMy8KWt7/OEHo654kLV8UJY6tn
wu4g8mkxofsAg3DRoROufTzS0udGrjLYHDC3FsFkkbCc6zKLKL6MfxZ/XgD2z3UlZFkGMVIMWY3t
j317MiwhnC6HJeYsrfsI8icyIHOeBy6Tkau5Bcepij1JzSlRv+3OBTvm7yP8BM+/BazEK+CaL0qw
anKLxbkkXNK/3j8CHpVxD1UkgxOgXAQaPNG1AufQzCV4rEj2kO2qYgLKdQdAHUyQbWRZiP8Dtq9w
a/Aq4y33OFkQw01dGlENygGeczAKBLlKqDt+oSFfYGX1HeZfqbOsH1VJXpQyuZWXhxjAljSZNyFL
L1nM+y22jswCK2l/u6Coq5UjT3Nv2a7dafGoq1/YzoJRIpe9z05UObL6oaIB9Vh9sc07CaJSI7hl
m/8mpBpX5WH8kw+Fy+iScF4sBL4VgSiygORa/HaC3SPnonNDs+VFSmlGuVH7iaYTzjeMVwfXC/HO
K01Ni4LUydKdwVpmLq9nmirFm6Nh8jpJjicqB1Ie489LAOaV3sJfft5DdestxYxVSAPzwU/9LHpW
MRQIzw9psru6l3020Z5Q7MzEPn8QFFtIHBPYxZG41l9P0LHMMD5ELU5iOSV+GGKSnahN2JnD2B/4
VslEpuZEo3WVL00/kxuERdUWa5RhaLP+JlCfi0Am55rXj20ezdwvhAknsSACzfO94vRto/V+Id2N
1LR1lFCpqEzVwfVVq09rUSEupsuLdAoQaJYXS9fiFfdgEsaVa9DURxaAap39oeFjKq6E0jmWwAZe
pBJ3/qRe88Ko4SFG+gxugXjyoTZEbIOmpoxAB0p4A3n6KO1o3YPIe/R8yAeA/rho741varmTMr4N
XPXP0Itv80NBGhbxD5BGDxt0Q3g1QsF0evxna/RI4vx5XOvAoFHz7xzoOT6keo1gGuuv9tWe/onw
j8hj1i5rmIapFOpm6Vh92ghdRydXS1EzNsg8nnuXJfWKvoZIs8dBMpMZXrQNq9tY3HO1bEQJaEKz
aPsZnz0OItIXyyxbhNU79wTvgqL+qsfq9pkpHc4YfVGyQPt6JdNEINPEUZ5KW4vqzdPPDQDKPqVc
ySscuimYJxZpV2QeHyocv0sRWnN+ilHyF+t5dHVsct+2aEBWfmT5mcNF3xqBpDCByLd+nDLaLcd4
NGZuXOHxqRcQQeW89IYpl9oM0/p2zLGkMttOwItASi+dLp7Xa+vrYYdgW0xssmgr+8A78xGcHlo8
CPqNVv6NjtqT9Ckk2S+o32a7jliiDkE0WNKlhAn/vHBVIgENVs8ddMLqWq5OnqijhLSzbVp6ViOL
nqou5Ro8aNC2YQPxlGb2VmtibjNyGIVKXZsmkzHoSD+6We/QlgRfWI9rgRJcN57k02EBcUNt0j8g
THbISR0qKrpXA+YuwKn4NkrXiVdfkgkmIdTxwmZjPGmNyBe52wLkRn/rY3dAhJLOepOp/NJ9kUTO
i7RnX9KEao1Pryao3FYbyJQ4Saja75ZLlo6xpEdDHV6IY8KpltFH1w2GcS5r/qL42goe/mnQNbFa
l+3q9+zSkpoKI4PPK6KhLhHyRFo8Ghf7UpByVFAPYtKUOqtF0qK4PHGdg2nv18rd14wItjJTbRnv
3VHlQ7TokRQbC6V8TViJietRtQYtEb/O0ga+8qFKHd+6LGBqk6nMaw7Gtc65Jn46hYH3gL8AsQ4U
/qxllM5fnp0diuxeTrWmPJgzM5Bg4iCky7EX/5OzXkrWN/bkHFB8xFOAn9PJb6XW4r4fOttHJBa1
mqIB/ab6grT9Y5Z53kQhG1joI7zV0/vqAjGDAv0JymuNbdvipGsiDPvDmM3zDRMQwhb6EbjnkQbS
qostQp8LXB5nAlzKBfVlN3VGirrNMUQUEZREteCPCrldJQ3UusJrsWFQ6RGE2mDEU+LS9kdn1+7I
Ol+qxgsRyHmBpSq5nm1px6h7dTb1aDFSDn25nCleEA/+dVE0vzU8eC5rW4v8b1+jU0uPVqgcqGrh
rLqZ39TJY3ySLsLqcIZoUjE8InwxWrQV3GbA9fldl0ibsL/Y1l27DYO6qHQI6Iba4GQFQo2hkwXq
8hpSa9+HHJJPlWjmlkCf4rjcq3Y21zc0005fmj1ywJjF3xV0QlsBX+Y0Y/ZdUvZkc96SC+pOmk6O
3qQpiRdPr19VPnINUy+QLfGDusmbkNCJdJgDgZBTkfFBnlRspVEjp0lJ9EjtItjdi6ALyO1uTpS3
or+lwoXhEg0zY7iZjO7qGXzph57Xr1fWOV2hk/UhrAOSUo27zUejX+wQNTgU7Gfm2VZK/Zk9LcFj
itTO4oIgZlKXirsPpUIz5GMKcE/nGzyNF3mcICh+jJ0WknNVQr+sixADas48bR0adEWB9qy2UWPJ
4nZ9GE4oTdCSsXGpIK47YsFkXp7Hfs6NxQiZt0tPyFNMWY2Tj4t4o6mRP4gBmtUEZnAmgUSvG2oL
VVeDr52q+hQNyGbQZ5/EX2Y7BADM0ssF4t+9ewhJ1hiHYuhNJtQQJuQoADMLmiyGhPjEqCSmtRkP
bZlEqBpn/G1VUrA1oO7+5tGgy4fQ8Aya7AoNYrK7zatJ5EZPDeDrQ8W+OK2RDsEqo9znSFvhaNMz
IN9AYGiAF1w3PP7jYSVWzR3lqwl7kwz2aqPug4JS6yN50HuOivGSjjijSSF0pyb/RfDoO9Dqy60o
KM+eW6rpKzXyx/GUl+7+E9zfA3074a12G4MXbGdAvwn3xeI4e/XW7eKChrl1zps+ROtgE9QVzkxK
gv/APOTYmw7Cr8IHqCe08WssnRSmhQ4Nb3Q18LAyIbFyDbYWUJbFiHIAWV/wNeOk+/T0AuBqCn1R
e+uF2mhjJ2qFaMaJAnNd0iOMp+sw0hU92K+v9W8j+Bxz2AGaqgBZISJIkrxM4QWphEdlyWSfxPkO
HQVjC/bvTsISpIV8Yrsd/LptpHDEOEupHu3ZI4AGORZx4ShnfyIBCGSOIjIx5TPGlPpcyNd6HyfB
C57G+BZfSWwnDTBAb7l8dzmqkXxCcXUbCaC7lkR4BHSE2oAhk33X5P3xovVfbbwpv4xmiX2EylEA
IHPSBJ+KdAgQbUesD71cMcSYFdRB/Y651vpfVy1zwPoC78/RU15HFntDORnULwlzNl7AnaAiKARt
hAM2Svtp77QWQ9yOTLoICP7gCKqw1iKpwFazvfhr11e08D5GXwCiOAI/hDbdY2pW+xLsSRxX2ql3
rnLmE87rVFqtEJSeeJ1lGkNoL9+7V+FAVjJVWZATCcfUZoIiVdyjdyJHzhVtHiF4xnvFUV9opqaq
c3UKk7WG36T4ux0zojKgrORPub8lFBL1jfXgXyfJ0wNrU8N7d9ubDB9yNhJ2gNEylPOK5HNXbmaA
KvIR9pM6N9ZKQPcwS6lk35XG0VOQdX6meeV8ruyjltpJ0YMXT5X+ymLiBHkISeLzzU/mVr0gmLC0
wCS2SZJkJY1rZ9fYXpG5vsEYiYfC1neqe7ih5xsjLJWiEY47r7T7VQRV9ZyssrzXfm/uS7+BxuaI
x6fmlQng9SHRFj/+47av+QchW7dnyjjfYGHA8Q3Rtt8cSX0t0PkGqiTPk/4zFI57QfwWM7LL2TSM
/Dgx+rxXSWgMJgrP+fPFdQBzLJpA0dko+XmJbL3BZ8AMPjZxw2EhRqT6epsSETFIDQRrpQRs0yGj
ezTfwCLqTFMMl+qAmP5WADDrofwetppZ7bd0BwNLHtgy0Q302P6GcMRV1ZZaGsnT/s05bzt3dRx8
0dgZjOR0MJHN3Q/skbGyyQpotdjlysQGbhoCVFHBTPXQJY/eNw2a9+2VyKFgU0WDr0+q5esfVIaK
rV+xo0Im8qhYS8+tsgJVBV+7Z3q1eV8O6hSkGu0vMfMnT8D1g8pUoOszaBRzMZlP9Yn+FUSOMVxN
/0bzDbmi9pSHTffHLB5og2jyOdnKNxtHbowtloIS+SjBgkH14mOp2CvQVEhFP/wPBA4jzjtssiUm
VrsGpKr1m6oEbboKdgCFpDmrdhSb0DxmxafaEpdtq2urkG9a8X32eFV8z6BqOrz1vAUzIoCybhvg
uHBioYbS+hFLzDgMmfvvL5SNGljRoHr24CGbaaTRsKXpwXZQADnaA37k/sp4vJ+cGVWfknojk2BM
jM0ugKVVRVM4mRq+YJQFsqhIQwf6c7NuAZOLptCk7chrlgkeEuIcN9j6O2GbaQvri+KileHP9kPp
o2ilWyzpZdZf3UtAeg5K6vaA5HUWUWYhhjd3KlLy6VIWWufB7uutdTGalvv4s/kCWoXz+jTiITtP
OikOoQUiBh3rXpdv7Hjpqlc4GwkKNSs3cK1Cv2uDnHkpWzrTWV9Taa6rGdW6xeUfihf2pQCT328f
3F3gOoR/+IF8pbpL/jc+lguOWbQ078gOnuZgA3NaYHXpIxzCKWTAumVQPFB4ARiiwE0nxHuwPNxX
k9vN7JYXF5hDgHjcrW1laDHlyXAyXVN1Q+5GFJn0zg5k0zL0tvToQe/ILAPNUH7vQ23rp4iRrFxh
ThN5L6iS/5dt4zzS17ZtxsEERMW21lwnwLlji6aqvpPGoOJpGFTjFV5ghRzzliKCy4PrPmpEDNuZ
5//m7yEk1VRDFmD1EKVrnv3BWLKwsFjGvi1ZGj5GFubTfIv2UmVXrNBDPtmdEVDB1up11ud3XdUY
30R+tSqa5nS/JWi5gLdD7T5iCm0cgV35RWgN8BKFkGj3qY1TTuxRVxB37IXwc9jiemt5nle5fmlo
oF6a2U+6iIWSpr/1it0gakEHU3bAuCglxUOJuua6q+FpGkfayW2XWbKxbmGciDErSmphLYO7BXON
pObbx2KhCb6X0glMLCCJ6tqpdNFVwU69lLig3tkmvoTn8i4It6TmMrmqK7+qSta1ZL3zSBto1U8Z
Xm6vuhZTmZSDjh0SFmKAREdn1NyMZouUfLBc1/KRxSM98Jr4mi6DlZGlRBtlppyvoB5xYxlDrXTx
+fIeGcgIKgIex1gHwTb+cW7OAsXApk7XxBP/QTlSW6JBjNDPzQZJ0GlN0kaq59JNkLL6SQpYB+mf
VupVNfaOzRZV9B1vTbzDiIAR7oeKLo2Co+x0wpZuz8EIVWs5NG6YnggKd6HcaT7YaGcAR6oMSGlr
x6zJxqMKUjn8noXkJGPJHGeZrdTRN+2gMSWRX0XOztgSjYlYkA5UgJfcbkzq1jr6bOrlTs3wLN72
nSCWx2aGVGHv7nAGrFC3pJEpeD9OdivpKUTaDUdeaVTu2itNa9DwWv83Z3JgG8zqPOHLRZ8Iz5AA
LZFqa3WRim2wwom2XM7iZZvJoo1i0maM4j7mVlyJqiyiqtKFaBC2A2IYC7ARk6EVTs/mCCTNxR1Y
hbQSCvf2UbEIceUrA9tbxy0V6Hxovja6TmSKPipojvNvsCphYttswB0fglewm2JvmAmORugPsG3o
rfc8CREqGTJQY/GGWweqwfMzAiD9U/BZ1TzJDBeuirfIQ2xrus+2sjpgmHlOFJD4Wx3/RlU+arXG
XSKZCsP9YGqf/DkhyKhNxMfiU1QZugyHhkJzLzT+lLM8JG/+Zg527LTyJg08CdmeE7ZT4OBv+AxS
Y5WkPAF0DDWCi6PAj8F5FyZ3+76tNFU76cO4sL4j0kYkxL2XYiLDCoSZS4ZxSjNyJpHqeSoJ+Jtg
0mDHQbder1Q6Wt3P3PogxdSvkqKh2iZZJlJLBOvEtSLIJgyWp0USbnCY/vMf/vV8GsoTJHRgFRtg
0P6ILWyOAQqL2G1nkBtXXUOgZClEW/vOgGl4EtP3qbygW8w0hsejETKZNoVfbpvipoKUB1VzOggA
UrvgInPWka7mUYO8wwKkjjRWwixrvrr/n0yCFtU7ixrKMjSiUrqArqo4WnIZ+UqAgvowIQqWA311
u4dXYXJi5Zzni584fcZGlu7ANHpMVwIiEyyRpLbZp7rNpvKl/iqqxACF/pMERl72Sd6b7rE3caJS
eR4uB6fN6AZ7WeA2yADObWSu/eK18dg2Hp0XnSx3yKR+1HEH1DZw/MpgVFQ/bt46WIwrJ99rGX/1
tUeoONST1fkoZL4idk+yX5EY2iiq3FgvZ9DgsHvAC8qmOcTDaaCziKaTwwl910wdOj1VDbKtRKQs
sLx+MKFGzVFosWw/H/cr/BBQh6BQMn5p84/7PmQtDBb7NmAcC43B2kO9j1fsSABwjLX1bB2uM6o+
hA26nmDvH3povF4DwpXoSBukvsItHx+eDghLUD7A5KJhWoFGDMwOY018CHkouee8MIcOBYjgZwQc
LDBQmF0EcWY+3fFrOFEv2uDjS7pW62kgicbD/0H0Z/LJYJa9G5z8Pqe+KPDe0vf7Y+k7leS9yaVy
VvcOSL00/XJf20DAm372GrKbtWLr2Bg17+UuAUsliG9kvsq5VfeDdKjuEI6aoAfOIbpZpCe4F8NZ
jQJyhJvYICkLsyRWaolfqTtol03VP6ye4vVqCI14iEGF09GI42+Gfmj9j5B8wLgBYjs/9To2rxPR
QZxytQv5ZIaIFC43fdcrCmWnuoCQe82SXflRmeT33ghDiBaPkgm0ueK+iD59tF5Xy6yGWGEh9sW6
s3EJ9CyvYLi0Yhi6wH+PZMzckTW/c9icCTjSpHq3bbWTrO9xI8cAuc0OakDvys4ignpiLNeVxsmy
nhvJDZeNDIuKSvJjgnuQemNJRJzQbUBox3UTcN8c55XUGKtldVwGt9eTTSyuoKH/J7XXxuY6ztk3
EK2MDjOvuAn/qit3HnzBYqSlwPOcf9F6psmAQzPL/y/AXvGrJR+XAdyY9OlUF8xFqfEnt+F0/1Ti
Tb/1LGVq5PTFvxOvsPhMQt3l4e1I9SkL6Y/UNqdMLPHJZSNuOoEkZLz2Z7yKSdVlOfSdtpM8OF8/
f+400ppWjfGDQIZ+g/BQ/csEx99pI25P7niZp208E7hysSGiT8/ukImEP1lgIj+6ua6zOFr6grn7
IY6zZMF1kMosUJI6aMSUzajORBmY6HuMY5bBAIfPVINMl6ktI857Ll7uWqWP16d+oNRY9Q7bLWUW
8TzSMtREcl82hNQD7ARAspdfjaNMfjC3aKnkXg+/BhvVAUAas2/oY3mSh1P8OgCh/7vOh8AQDOOt
bZDBGDnNZj5ntk3Ss8WWCrxad0g+vTNK7oOWmZhKN6OzREOwmpSrHx7I5BKOF8vd+KEpNxu/PlKy
MhprU5MdqxE32J45CV20yiG/R14bcwRA+DYB0N8yjz5lxi1Ij+8ONPBnBGgKEo/Ga78AUMCw0t8e
q8JyUIJcs+QUpctzRQbpoqubXQptifsuVqhc6OwWFIEkJ4MGxKvXb3qM2+4/laSiSL82vddRdKKZ
88jg4gKFnh+wQJULwCJHEr1JdVJ1Zz2D/vuIHS/wSwrEo/maPSGmE7gGkSevW+iTr01Yr0GGgVIA
2dYOjxUk33FxTAyUyUdxdKC9tkBGF6vLiE5T/do/lToSqxft6nIOm6ukY53Lr+Hccq6mlumSOyja
0MEsDD0IFXDH34a3Y60h6zCjhFkR7jlae+Oa9DqJciYX63YkJvk8EoUQWXVnqoCr99rWzlH9fNKb
m61GNbHgeVzvrkKPnOsRblVe+1JaALt7ATDt5EKrVNwYETthdclxGO9pi+1XobtuVUlRdlj/siL0
IaVGT6Omg7cqwXEzEC66cjj/+JVh0WxqbQC5Bo+81QYPK2NKgLCY4mKHjI1oUKsQPbGodAuMKdn5
5KqNCyOv8Vs8vDseLLnFnvCTIgpbbhJNdUD265SjeVTdCwjq8JxnjMUPAK8rIR+czf1iZj0Ff05v
sXuGyaiT1ygwnIA5LLy4bl7UnE+V+dzQYrJpRBVSp+Fr1oHl8AvovI8QpPi/w88LWgwVrl65ALot
zABOA5POQ/JqgHKMRHrj5I7Yk8Yaa1IOcLc99kqWQomLiC5IVHxFVwhYo3Ld00P6cFW2BBii9Sva
TR62dQZi/l+CqWWo5zKhEfA8aA8Zs7nlzqm/m0i8kMkBlFx667Gl3tZaTIQ7kUmslJRRQFDZRdml
8OGN5EPcdqcmpDqZU2RXS+/tpcqOQjudfNJPbvR4ubOlMIuzRbAFVXu8TcPTP6qOarpPQVgUpN1o
5iCdXRmpQCNgvRbFtfsP3bdTX+EyhJvjzKgm5FHrAwFrgEwPz0RLXfmKKf6Nh43hnGmZRoR9FUvM
kk2eCaong+X9IB2ZYhRglc9+C/s3ZzQ9ps5vMjgezw1RkEKZ5xfgWtwZ063qH7dDyBH7kktxbLhh
Nv8Fx42dEzniUTobcPYk+Ox1PS/efmARcPq4xl28b3dYKSrrN3/etEWaOOXwVcaTinY94+UXgGoY
WZaB8R0Qal/UvaEGVCCiO7jTRa6owbrpkizuLeWK5/s1jghOhypj6zHgjCWDvjYTDrTjE+rt2mIH
MHrKKdi86sbx3aXdLeiONCp87PBwY3SzdTl5jRNKm1h65k0G2U0i+sGylEboUe7hrYvwMX3MOreT
UIrljJxViBtQSePJYgPgabzcKYeQSQyz3GCFjiWgj7y3saHNNIiVhgSkfJWbu5XldH6eTlZIe3ER
tw3llIKqWztK1eUsr0ya2LFSaqPK+sWcFoC7afyaq5g7yu4QALM3QHTMsmMNWwB4o1bYrRMmmMDi
73z/IEOdrXnB/MTOfrW58ArNiqXqanz+jwUjmvhm5rtiRCE9tdb+BMCSif+whEyLTrwVzsekQqFh
brgm0akbu2/h5TOQCngU+IXUu0lIkwGjSZsK4jWHo38cI1uYtEgp36ZuaAsYXEUKd4R7NKgYokhu
rBGrOXqHJkEYZdnNFwsWBgjw6P4VIFVAU/6jBg3XBtTk9Tym5fAT+tQWK3KvW/KOX49XhME2FgDi
Xg6QifK6LYs5qz+mooyfc+IG9xy6wTqWXZLY2xCsIVrjq3IIO7Efo1KCA4Kh/Qw1VYCw8K5uXjFo
v4RegqPjKyxgfAjoygP9nvd9IIZPX9PJPNVX+odwUsMpIZxAVZxEeeGytV2skZl4c3j7PiKTqsFf
c+2TxwtsnYXJcTAaaaWkRSXuan1/f3Y6NVhxnOLyK/gxSXsmlWnChJAppcd9KvHeFLO8ClOdKYsN
DHmKoOhvUvDZXB646L9ORT/sD2lsR/f/gIZ9ukj/iXpi1KgsjCoL/e9p9BC5pwcTGb9R4BwqfwCk
qXQv4Ba8dOXCYiGR5noDAlp7Wa8Xv56gYhf+NkiXLHu7juA0b0Rrxh5qQVgwxuOTNXyftLFBrxh/
Z/e/esbVMOt9sSr6/8sO2Wk103xc1A+3k5P+5sguSk4BHL+uQTyoA8iNjw9PGFlckuVVW9EYQQuo
YjjDEL3A6JQdjMzX/bw44+5COiB1iXhR1kQhl2Jmn37j8YULa1xinDo5NhoZus8fDJcjfTgQRRzK
UlcvouAXEhtLYo/QHu5oNk94HErR5OTD5JuCZeolWXCxfT6ulLuriFNSnCDuSKx6gMHDgtSzEnZ4
OgU4pMiA4u5zHGkDZPNKO95uTy71z2ueUVMDYoqT7pxjj3sU+Nq87Kv7ks+34ADU2+T13pAI06I1
uvN5oGE3H8puZSFhKvvjjMsbxvXbga+xNATJ6mIQNm97BW5vevXGvv3HYF4LR32I//52ziBVpmz0
84N2GU2TRTUaiJ10/EkOgQA/BMovLEVMSihRphqHY2nQ48VE+wIp72yCnHWAyl4/RM5ddrlI1Lma
dJp9VYzg7JLYr2DwGtwQcwJpHt5HYbpFnOQY0UHIO0QmVWhu2AJf0yo4oafNEvmSAh2cWE8YEEOz
K7T3ag/xRBO0nFOL9Fd81WycJpLrnWd2ShjrNRALoVf8BJjJo2P8WYNKvbA+qka31qEbgqLWUIV7
vlSBCKIjPOwtx3ebGRaMXesRxNzaL0JPpI2Z1SH1gHm4OnI2tI9JJfpfQT9b1MCsrnqBOwR8z4km
NKLDuNPCTj3pqnVPN6Wkbpy++X9RGPKIcn8u7nKy+Xfg5yASE/CbfP9688blHSVrdBu9q1cVUKiD
7Yq1UwicTQEa/pmh1lF68p1miyiOe+b2aHAUiuBUBwknZRN+7SObBJBcBAAKRbGzpJs4mikte//K
mI5uc2kIN6fhxv0bCfr+OXS0ecaq2e9Kt56/mfmd5egs+rIJuULvnHoDS4fc2+cBgFVZSQNpQLf+
o5La0ctkMw1ioleNAbDI+CBO30r6/c185KenduZ5yDZTm58poQnIsSPMgHhm8PshxTwkiOBSIHNe
gyGCD7ODAkEu8/EyF+jcFobB1O8gbmRcrTOwpG1C8pwWIMf1nqjODyGe1oY5v4tXI1x27RDeoFqM
UeZe3nos+K8Wc6eq4CTYx7Snl7RAJL1jJk4P4jbait1lCrfXqtrvbn9DX2s9PLH7ktfq2zpMte2V
VZ5x394Zt7jrksWHQS1tW3tZqYqVW+CHnJg/SoiAmbr8N5cdM8eaYtuXeLc9cYLOccklS63Z0NmU
wIqCZuANknRXFwB5Z33jws81vw58l+fWuu4ZxXML9nf8qWTWRJBhNxZHssjPFbTfm6tRgNZ+909J
VfSEHP7Owljhc6Oc1pqrGszNzX4g3GQN4jjTL18VH874gvsOK3OBnXZyZctg9IJZ9TvM+xUdSj77
K+yTSer8CetDF0+15RwkcRn7XWOs4R2KgyNKC/fBkgij6cKQgXlbXYpQrdV2cyL7TpQCjfxrd4Kx
tVYIR4FjflBzkRF7/gq+hZAWPHq8oztwN0VFdCsR8s/jHaqqPBD0YJGX6hxRWEkRVj/zGsY4dfnJ
HOcej9kD59nnSmtfKoMvWSVxtTLfbXNBOVCZLlbucmtEIDftHSv8bfMugOYI3Rl/RI0d8p4E2dkp
Z7odSk8YBqssmUBYLWou5VoyTkrsFtNfxzw7ACdQmQ3N3T1R01Tm/B4jaZzFzCg+sMLsvUUPo+l0
sCqUh5NdLrCwN0nk+8TkEnm6MQjHzGnDJTCjb0JrfvjYQtIVEZ53sN9XEWX8TWf15ypx4LoB4qRI
9rUsNA5UyhSwoc/eCkrY0kE3YDv1NWsmrAj444zkTRhvKc1n+7TNJbR6shMv5iLhz+JlLFXwtWGE
AIcy3sMeSWPPMaiDJwzy0CsPjY20EKNiHxRBQy+EZGxTFjliaBZ9915IhpZ6hGYvlTqMtMN2rDz8
y8zCo8jAGNBgORvNB/o8MOTSJwV723gvLeE27RIeV0i1dhzO/OHkiFarKE0z/YmXEBfZQ495IBBl
+9HiN6CGtKtdu9EqkIb9t5GukR0JTsX11JvpvY5EXlOifeViEGA2TQzlv5GSuMaHc/P9q9wd/yZ8
shWMErXBOdxBnqU7GRg2s5CFR8SHN3yOaCijE2I3gknceLQS7E+aYZ9nZP+Ha2PyQN5g+gOu0guu
zRrhxoOgnUn8AD+4AewUMQ0Z4f/t5QlHQVjUL/jZM/iV0HzKJuOI7EmjydJ+qqArUpmmAIv8ud06
Vge8HtpOxuX5vh0FlfOf2Gb32L3MC7rkdeSWPZfFtoktz7hy+eXKD3EshiSNHllGzDDf9ncz5OEi
tSwuxMqWFFJ3NwL1Cs0Sm/TMuy1FuTJlsCMamJZbnNvlkCUGM8lNH+VXotF6lgN2x0B5egXseiNh
RB+MRMyhXlRf0vl6Bz73UYu8N1ZYnnu6b0YMmhDsDAx7ZEGhz8TIBGtRABmr0avfBeAIWqUAMKaJ
i/HvxOAvKB776GpA3Em3yM1tRrhrz1Esz4z/CFeX4tX2v7CU6ndd9jMFAtawx5hLnBG8y6xJqNnq
prFXKxX/KApHT8wtp695UQ/MEpxCnJFsqpd+j2MQT1ravZNEgmjClJioLZo6d9rb+LGkirwP4Glp
kxMkypVpSlJcCheWOphyB6ZuVMet/Ehfau5lKY7OO3MNI5e2tDYbdvR+rCq8nUFjToLtiz3yGUFx
c21F/u0iR1VXprcEKfKmDlwNFKXdCQvjFDsYB7A0+kMnjxi6O05jx089dcXpxnm0lrXrAdi53fqP
rn+EnDnrhYPIppPVaHKSGrAml09wDoIcpha9/f7C/ZBc1GSVhK6zLLRVawdty8ZjTttuHVRU/ek0
8ARUN4b/Z0J3p20zVmaVga6qlndgAPfb0jHvtQk4sM8Jkl/yRxD12DpIO9BGKMuaHYJerQQusbMY
ohOsWFAeohjvJ/dpMtHd39hgxzPIg4X1E5zupz4NNEzWGoeWl3dN5qU5vq82HfDAnjP5nGvH5rTo
4Wf1NlnxBsDZVlvPWZjLh/k5CaWqbt1knQPWKB3+U7te2V1k+pkbVU2kT9RbuVUL6U7N4D6TMSMs
acW6QLu+BSl0AO+w6WJoPdVl79ICqeaNmVFZejuXPAcdHhnxyUSOKnBuRRutIP9ct4qtZ8tQlEGw
rpaO2t5bjzSUUxm/qtwBlO1Do4UKpeyfplt99t1eFHBrAC3EW0I2fzf66G/4OoOb2gsxv0vBYjNe
ITnJWTeFjtfX0NicFXty+xB1yN3UNrT1rCGa8ZxUcJbARt8aS2MwhtBcD2Kw7h/EwqExDboeXjrn
riBLtPxVMDSpLbls6Xh1JnU5izrVxmurWCzN4XzrXq13RHSFixoO06OMzvLMSbuW+QNrkNG8a/rc
QIIsSF5Ggsly06Yfm/FAyXpV6OBfRPBDyFxXE61cNbENNqEBMmboXaJR8z94thSfz0kzSHBYGOj/
58UuGgWBrgaDEW2LqcEMN/TdfQ2b0B7pu0zk36Uhkb5vdlVdJHF4l6rAv+HnQj2cSadfEt41R6LP
112IVb3j0eVt1gZqPUJywTx53WteShY/P/1071tAdyVrmk2ArJIVQjaJBnKTH3psBeJE3KI3FGab
oMUonorx9sAAsLQOknxBuxDcFnNM+no64NZlUmRhsESFl2VG+zLlLP1eSvH87U/2oJgqF1O2B75K
VFBoJkrduKdS+twlAXeutY+tQzwzLRxSOjq21hvudpSqaIsWdxrpxYRxlHyY1po8r8bRXk6GBJQM
W1Ug0jlTMoHpNDI9dK02w6BKVM/SnblBusKV0DlKsAl6oerPIRsdbzOItEUrcFy76JZrCStukk0m
ncZvOGc7dXlAzgwLQd9a9cOtcHeHnpthiS1NEPMABikuR8ZmicfhYKxKZVJh9FTQHBLPYltzPxC9
aVMNvfXNJy2xPNDmBILY9dYZKm/Zx9M7wVGQ1Ccb2Ly6/KKZCKH10JrgkwtnSSn18mOZMOqFWv5S
LADUIJWv3DbSfuzPXcmpRcx3JkzFtiKLdXtczCb1PwbglWj3/ILiSKYnVF5EMLK6i8WCC8QaeTwe
m+PjNY3YocUfC9Wj3+S7u5t+xFh0oHYzQn6ZBzcseA3YSBPQFVozYHYY2szND6mc8SEThRARe4xF
e+dxCB15goQ1g4M1ssu5Vayww4UHKZd4J17nOK7FL6fm6Kh7O0n+Set4TZQPTCQ4p7+XNgF1mAf4
Xh3GuGeV7vdvfUu7Ca+aIM4maGbOkMmtYeCPvGAdhbadco7GG66gYh8nRJM/UyJaWKYNEqHVsHij
4lCZjXDySSUHn0cXm1+kDGc2MbzxwYzJE9CL5AK2DyK2eIj3HxRt5uopUuL6IbnF4Zxju7mF8SSJ
f/ISpdgvDcDv52gEasWRPiNhsVM/hYiR7pFT7CObA1qxsgHYNUZNjvhYPVbKjMMa11AzBu9isfYo
f20A9f3OpvtTTIeCyp9I42lXOjOANJC0g0DRxjxcAZgn5Nfvl4osLmyC6x5fpMumJKTUayGeO0gt
FWEJQiMUDMzU3ivT3Sfrr7iWbsuEnQF+mPot+NxEqhzY3BY5/XWfkXpsxWDQiKpJS7fVUR/V2Njt
dt0vJWIo7thZEEgdamdfBK0HJHNDkdgOHmNCN8r4cEaAXXTKSaRUoTzrVpBe2JFaSvpop/bC9h8Q
ZMnTrjQRb7whSv5NrbH0rz8AMFvOysVcrANeUzhbZwQXuKnenv4Xl7UBmpHg6IMcxrm3BZOih92e
mfhNQIiuZdzp3Q9Aur+odv5qnAElAE0jzFhIUP25gQ1FRy1hfGiN88kSAktcxNE2fzleFwGBiLF2
VdVcT1AirHWi00vO+kbX91VYJtrMf0eZkATXhjUM5+xvqrYpUJz1H7PTRwxUfNA+vI7PNe59iu4f
Hf3KqI2fMUIkMe8mXCxl3Q7hUkZXck0zcUwsyYhhsqTQf5FkOUHirYybFBdV0MllZGM6vXqK+CNM
lP9jOaptsYEJviBsKD+uKXu+YHJlwLf7gjzIdAQq0c71sbaXIV8eWi5bi7s03gjnAmxvENe1Qjrq
P9NCTaxRqoBpcEut9NUQeJCmxQRvG24v+BjAI13OiVfUDUWUZkdCgQFKf7l1piI/2ktxdfc7eFsR
LdMOWSmG5N8yeeVfkljrvx4GkgauHWuMl/TNpDaPlOKU5Mg340Y8soqTP6hLV4mQaUEUc1KW49RW
Wf++fhHN3spXC6mQrny8XkT2bfu383qObkjlk5C3rJHxl+KS8xSuTwn8X4pD8Djqcs7AwT1iq7+2
JkWY+Kdibw/wLI37Zr1SoJUemdqgYyHlHIoWGLUwAzVpEtRAoiIx2OWi3jb+QM32CkCdXFTTYaKp
3iQSGkeQu+/Y+HvQFi1YDZm83BFriv3KH50WsgScAlRKixGcKle1On5sNMFyYZdjZMQhCRTPtjrE
38N5bJ4g8olDEyilxHNHyNdQHIJmDMchGrwxT1CziHV5vxh8H7fKYiHkf2v7Guc7xD3u8R1RYsm5
Og7k9+eXsEt2VSrn5IRF0mkYt3SDWDbtlC7rNe8oWx2ptChg/PJ3xDoBtKpiFnN2C2khAe1Q6AKy
0QCoBD1TgB7PN1j+wvcNToHN0Wj/Mq3LwwMU4JeJM8uv9kW3w7Sbe92PslulEwEa5KkdVBrTrc45
Kb6l/6/yDptbdNpZPlTcxlDna1/pRF8O2UG8Qupgkilm3j2rVobcm+kuxWMRd6hzSk1S9DiUS/bS
j1NDPysBxFNwCzQTGopjv7yVFIybTa03NedjuwymnHqeQ4NpyvvEdcgybcYm6m3DcOb8ST+BDism
vLFuXkbEscY9mgc/7SWP4wTH6VFYCv2XGx3j5wZg83nm2703vXwJ3c/F9y8gK3N0mIILdxhY4cJQ
jDkTA2qFSiX3apd1R27hVRF8M0PAjYKuMgauAiTh4POkjsySG746wVQRpLa7pW3HK8nabq8q+t1s
061bgYwNi6UgROakGswegvorNdU9EDYLxV9YhW36xlSUehkyCZ8AEE2yYhA03rhkFg8KoaRXfpEV
+Fdq0TpmsSm/iO6+yMspiFKw+vzI7DuspSa5M1E3NcabaSK9fkqa0WseCN3cE4+aqzQqoks7OJuh
4bDuzWZ2yspbkP+1pv9MTZ1E5Xsnwx7GfnjZ3HAUqRggJcNSkgL9HNGaxkuBxLRyeuwB4gg9Fza1
YYfvVdApZhmdYakh3OwVzdUotuC4LfYhjotnhnXKSqH97q0bwzNOVx9eTRYKNKEsTvHTtAmBV4x0
5CoMzIkJPwO0AZSnBWqjPQQ7xNnoa1GoMoTYX5NqX2HKnq/7myT201XPkiHBqK2CenN3kZ9cpRdM
0lDKjgsN2iitywE3fPJO5s6PFI0vsaaYITck5v7cuQ/O/e/BQl8YbavamcHQmGHOosJqgYpiePG2
8Rl+umu7ZORqk6ht5XCfe8PxrHLsl8P5zZwQfxFH9G7FXnTtJZXjRDwVlstWmXw7N14oKc9EXttK
ebpqDXG0vhAPwvd+JME3jQd4B+CnxVnA88rST2upBrtC9RuZ0UmyIASPv1XB+ngccFQOkHw1PRIB
Auw2HeY5g3oi8haVlhfDyxnm6E66x7gIOBB70YNp/tNlSCRF13Qh/QpEVsGz412WqliXXeQrVCEI
En8nF9OJYaZY8KNF9YQZRI8m0aKxKp6NAiB/DfMMVqfgSFBrh30uMRX7WDCoUZvJnhFVbFsgZ7WC
vXyVpE+rRNacmd3mBhvXOqqRyBZ/6uRL9rlMlkEfmCChRjT4+d39fOGO5bXeJXs28eDWqkgygcJw
77nCHxLcZnCdR0qqmhLBowbDfOjQvQD0Kg68D3PZxfIYndTR8Bsa9RbMmCir8c81HosBxgXniZ8O
POnG9RLjt6lgfq4+9UWLGuS1q7bYf0yjiEAMx2Tn5IQBcr6+r4TP6tuM6kyMtFQY3SwQc/FC1I2U
vEXG25sR9AwYtM5BLIFTA+UrbFP/j3RGTrG2OxZEuFkFP/cs25RQCC/apSd9QFQfjdGhJRT1LdQ5
AZMqKrsNXeS+BLdEV9WXzlpuZuyPx61n3QdC4P7sv4zyPq1nbKXdoJdZQgckcfkWBb65/SucftSy
gu0TGrODVv9qg4upjiNHZumL44RLBC+QBfoOApTd1sra95lWzQW04rPwZ35BIXBM/xTAzBzvTki8
FZX/Z/58uMeXbuT8JCi3oVvnl+hzdE3ciibHncceXr2hOUmvqg1lBbIlcVbfuSxcVF2fkNi/OEiF
LypaJltlg3cyZJ1wiP096CVCoyG/0v/fNN7A7NPsZup2i9CSkiKo4ZW6vNz/zkJNvpqRa53WR4+s
HMeWEVBaNdaFGyRgq0ESq0o8pAusop8Dk+Mk6JQzqVxXUvtWZkuBTNUFFbLgdsFlWlfOu8SUJCB+
odtvBoyMu+LV5pRPRwtosm/JjgyABkWtBN/dErFuFsTV0WyGMe8LvNeiQvTC8PXDTYhG9njtXLgL
jjMuoCNbT0y7SC/ORSKCGkYN/ytf1KGUbHIOyoRJDSvh1aIclWdK+e+XY7daeu7RQZKjEkpF3zxt
FiyW4s1w6ZafGQNkfICzzjHmzmnlEq/vR9Zkm/FhfZtfMnr4NpQMvV6h8wH5iRghc4RFmvJQ19hA
rgIao2liRIG2OWiO13agpjI85Ed3gJWxhfIWdJzhJqiIAINTejed7QRrzC66r6N9CDLmWmdBKqD6
f7ix1h5a5YgxwQS8+wOWymIQ1AxAs3eDPdM2MgWwzPlfJy9ghzNWQqPsBaaNT4S51WZQSWDmrVZh
q5BV/dSSxUQzyM4zEmp82h9AgrRjhQtVSoPRq0467PQS7Ic/1OcUGRUsiBE3V+POnutxexprZJu2
AvdHUvwI8vng+89ArKhlDlttpaHO6Nzf3PeStEN4ZCea5QvrKAgXTIZk4fu7BwJ4DQq3z5wvgFNz
cFpiYcTrmHyQSbisHCgjn/fEvL8/rti1H0qX5AK6HY/O4J6JI7uqvDN7oyF6XjmAYNSBgwJTQtNg
vaZoyppao0Op4mmORahV8ebnvbkwvvd16DsAgEcsp5UPLXr2JRBWc8B6+5pAOVKhxvv0fyfiFWoF
GoPYTFrmNZnqL96euZy49mcfkfGqPNrv4JUQL0NpWrfJgDVldoO27hNm5hVOoByhc6wDFL01B9Nl
0rAU4ziWNU/yNPWEQbu6jjclG4XZ8ziU3j7jaVmam+C6xUZhWGBQg4/4HgllL95KJ5wA8J6d69nU
4Jd9krQCvGMrAhUyBdDJm14qIVZhPUHYxgcT7yubH2ACbu70C1nMvGdCsF9VWqhqt4dEmZnM7b1L
/tPs+al+RwFsbsrT6UBYJ0nt2MUPuRfxPIk4sXzEu00tOj9ePGE4yXbB496tsMP89+8c0PqBPLZN
u97WYdNFyYRGzEkkES1IhP7IkIWYGnO0dF/2Gi09Yxg0cjPxSFvnd5xeMeK1CWJtRatyU2fAxZv3
VclHlp7mWGyF9WtoaUh2Gc5Z5R8HfpsIZqlk7mRJNqNLnA778sLrbi/okjxUzddy63U2ammtojon
treFCtANzbiiNUZTiqp6+/LVpo97SLc/LMF69YyOnusW4iYFd5B7n69rV2zRQf2WaZa3u6G+qMRa
DdD2KkuLRTgtn5MmjtUrq2aDouNhCR7m1BqiVpcNl2b+ZXM5yrG2STdYeQ2nygmxdcU2PQT7yKVE
SS/+peJLy73tGoTdq9LOWjCENo4vaeaR4vu4SqME5fGj0WQvvkOD3nropRZtcL9O4vFWERoLx81X
SYGTd6ffOA0e5H/X/Vg3K0JNvernFbSfM+3ph/fp5Kok53+3qxq4yJGbHJ6ncPDu2ibPXX8QX4gr
DkS63ikTqv5aRQbxZsBP3RKj9hFsZAPdgwAvIld4qTxm4XV4QRsh1UB3gYupLPCKzRMwwzpcAe64
gVhGeiCwEHyg7CJ/ef/NZflPjrp80eH1OBdaeWlnnInUAFIne4jhG7Vivqx99nj/jm2kIEZZpZFj
vQ5l3qAlb7aoshDr5ves3rFnfxQ3WtqmVBqrwUfIZJKMLXb/d+ZQTeGUCJjLPr5s7kuACjhDF4kt
Lyso4bfg+YFA1I6/dql/ZgMP73xKszyXaX7ZPyNXflZR8i0Y1n48YpzaC9D9+BMb/mTlsXNdJqUa
BG8UJ793PWrn1LSM6KFipIu9E0wMdjkLuRKftj/VKq75AU9ksgsdINRNaTD8LnKjNlNyCGDbg/pH
4dSC+DUO+rg+Y6Nwrqip+WWZbjswkwssDZiRceQS5+tfbBh4nh56C5Masg9tvxmbAtlwKtKXePm2
QBUXd4MUG/mqRKevFf4cSiT58t4b0AYxyT11pJqoQXCQdnIqKHK+JlLO4Rp7UpvAMrERuSwljSYQ
VLab5WYwgsi930td6U/Y+D7FimWbZPv8cG9iYgjjisUiMebYPd11slLAqyOGnBo9EJrWZeCdZGGp
HNwd6PEzbJMLoIFAN/VRg4uTZYdIQdR9dbs9XjPW0qLrchgDxqv+eTfa3UD3K1mQRYfmXQX4+KIq
LtCLLwfZX9mis+Rut+MnrA/mE6mmyDoy1iBenOmPCRvnSXGjbLZTjlD4u8sh9Sq/k9HfBBgLZ8P5
W7OSK8UYVmw3LJIA+4QVAWspGFEq2T3ZV41Ydc/6zbNvr+yux/Z5uJyq2UomRts36JqFtvXtaXTt
r/GVbe24DGg23waJkyPD47I0yBESdmOJBP0vVsrK6ft87uwi4RPa9OagxvojTGnk+M/aCC/Jsooc
NBUpoNNM12w/hTOeG5d/qDcK3fJb6PWkUTqMLQsBFKwt19WGfZBIOj3AW7w5Y0a7HtwgRKQ5hXxV
a8vQAS9irvdGXMFKJiHoGe5HCUqS7SvNCucadrbXl1J/f0UcNs4CfKQlYW6XwdZI+y4jgtz196km
B8ozPYcfdDfe1Dd4HUErg9mQEmBx7KgxzpJmjAc2mhG2bXkLibgv9amCA/0UsHqE/uEu6s5he24N
vtSQ+Z/7byvcJjAYBKxJgITrCKoNUUejJEjhFMPNRSfc5LrA3nkDUJxiu/Fv2Dwa5i2pN406xyNw
9bhamS7mQsEvIblmgwLKPbiL29+wl8ixx+BU/V881Yajtp3KAn2bpBHRwKT6Eqk3FtDSQs1zQVm5
kr6B3qnj4mwlfr3vKvr4Q+FFyYUGUrSFKJVT1dNEqMNh9YNCiBQJ89pZnVyjfnxxl/0EbH0xsEy/
WaxbnoHkqK1K5D2PJJzmNQcNhddW8XsRp65bXhns59jy9laoUOzalJyI5r4bWcGT3oGtNeWBIXKK
dwWEeOxluuwjlvV9i59CkAgzcceWsxH9d5hiU394FiyBvqXQJ1pggONUabzwuYPkw9qsWOHThQg6
XxFp2cIi2PazgbMpvCcxzTYPw/9RV5EzdjkqEHtgc6Zb/uh+pYi7bXYRJpdLlgA4495TeaUHbL+V
YEH5kPicB/rZTg9ss9uVirL4+DeZRfLEoaqYfYpdxyXU2HZwVWIdciIELmShYew1M1X1vQARrLVo
fUenAtZthAzgswDfiKhkiQ4LGuHbMljrqXwmoLgFhtptsy7HjfYATQeJrb77EaEZQDE9IszUKIKR
JrztxOBNvD8iCe1VvtTjSYCKQo+HGSEZuvX1279NWiD+5ZNWnl22brq1vRKE084AQ/hWIBAxEeFd
ImSHGTN8+SPAhDQ7AVevfbZk0JnDnLh/3HPPpIyf2+XBQbu0RvHpex/nep054xIMJYi/VdA+OXc2
kQ1TL6/C2C3Vx/SsVS9NTqFlQDe5IYMHqb405y36YI4/E7xkeEO+l33WsqBWakXTYmykcxHn3fn6
TsWO4ZXovHBTgkw+NQdrdjRIhBZFx37Ls+YcImWezM04bk9AX8kAw3M11jra4yOWTfw9Hk6X9Rhh
qWHh8hc6bNPJlWRLiSt+XsTjo2FgbmJAo+sX0bQjk5lhhAUZlYNUmQTKOan4ZIHOXgFU7AcMNFaD
zpqVm8PoZlgZdg/BIO282AeTnegUT7FcbnaaHAyWRmuYTAGBNKXWVjFyqcm035Ln76+hUm4bU+G5
V+CYYro8xYxYNRdXj9KK2qNg14eKTOur/LiqG2FP1fiMrf8JvOGm/tN1y62HBfz8O2HKqCcSNxrW
vCIULmttVpF5PwiH139ihNzF9SgpdE9xfFINhNzW96KY1vEZTssdKiTKRqdZd5WWf+Q5LE/KEema
kOfCCrX+pCf6e7+jbD3vOuLKo7mxmKHdGsGRiFkj0y95zaRI8o5nUkH7EklMYI66Kn/M1G7hzfJ8
Y3B/dWgEQKLGuXooMhPMNB5MSz74y5iwWtZ1SrYk9M2PvwSVYJ9p2m8uyXDpNGBuRl8S1sdN7CaW
iG8fk3U/3vyz3/6pPEaw1GBhbHGexjMlFcCL6GmBnoMKOZqU4SkEGTd9kAzc57vQhIIKCmho3X5p
ZgJ2P8PKvTf3l5WdAo3IoPTRhPO17qXrUdvBoehzrxqLYxktKJBSIpCwQZKkVoI61IIoYO0CmQ31
aSN6wpphCoPwWyELiXSD7dvF0bPmrfTOnvlihdrBJQEVyZKs+BdoF7bjaiHdbCvqdzI/Ht0qq4B/
KS+1gzhqzjqL7TFOyf02Am9zdjf0kKZNBztf5HH/8M+RSFXaJ6V1+veObNxeuboVzfqn7xj4e1QR
fpUGOIAA1JqxEN91Q0lPJ/NMpwT0jof0RYCcFMSXUK3AoU5Q+tl1JMLiQSs82/0fmEcNAR/qyyDp
Dxi8/gO9Oa8EojHhOJXv7S7MYmFSbJ0yXxBgL016FrZDcBzc7Ec8jYKTokutA+UEd0Dku+Ae8mGv
hQuYHuuuVvNg7uJ40tDFSy0TDt4IK+Z6FCHMtgv5kCBy9ieVEl5mcB0++yA64llwEQSsKggQmNMN
gjSmB4ZKrLQ7X8QCNtWcotKgxqAIPnemmK/2hUZJ2jfGGpwM6aOISZWiHJzExtjbrtgdLM11tgP1
H48cJ86TTRXjfgOoC/lOx4XM0bECnhKEs6W/wl0/aMB4aEhBz4B4EvlORhPAOEYj93Pq0JaxWLJ6
aH5WwDPHEEbAsX+XOdRCwqXavUd+Aje7jX9PeXbNemlvrpv2FWwN0IwRmFTRUQdp5BEiOcQJU01e
33pm5jzp70dZKTY//39sO7hdSa3H/txooXWALF4oSqV5RwEl1JW1Zj34b6lFXCuA3xHZCtAiLW8H
JWmBE/mbNqR8LpfjDeY5x+Kxw6hlA9Obv0/MwxLYCzTza1SVz1tCxPWwz4YG8zSTAU7xzyCejIgU
eZU6SuXQ4IF3qK6+eHqZMAPLnWtA9blBFbB27IIbnDItqAHqlClSJ6aQHIqZf25auZkwhIssuNGK
MosT43ZlijwRqh88qehNVvlbv6i5zSEkPx6suc9jtc4/rJzCrv91UX56/ByGf5eJd90Z+8lEiKGb
RsJAmEyIZIU8sfN7+uW24qD6qT7PyYc7mFnXyj91XyohXD8CGbxanXCnoEny14uneIlWOSSExDfF
vd8oYKvHC5z9c3H0awpT/T+3ZtEmQE8JwE7lZN97AZGcqy31YPk/7KvGu2Ri4T3skqwMerxF5kYV
T/DHShDI/Eb2t9+KNtRsheU0Ic7b3U/dukba0I6S1YYglahthr5LhHVC38YpZmqup+0DiEGPJieX
0ZMwbBTLWfQk/0IFw24RgwZJrBioSjFf7Kydy4zwem9wAx8AqK9VYsUatlMMqizmgPxzi3f+PnjK
r80jcDJNJMuoP+BHPCudoFNRSA8L5SqQ3La+fP2hoPMCCPPLQv/SkIc2zo+0F9y6nLMj+JM70l9e
tubG8e/oslEQHfGl7Z1yggRBchOycuntRYc+NYiT4WA1/07gW6wQkXnblEMRcvXunEZ4EOmcBttd
OzTb7Fe8PKRt9Q5bbV9AcTbCwFDDdmPGJr82e0a9TrSgK2ZAarX9EH+Uykn3/bkayyo70aEHoN3M
V55QRRiZk4YkebLiwgcFFi8Nxq1PMUXWoFV0IJ7JWD1fN73CeNX8tZkrM581cleTP0nswAd4m4pi
ULDKU4VZd9RNTj6KIr34g1OGRn/EX8KWwqUgpojCt3DFlW/jKCFxccSfNicN3N485n4A0yWKJS8g
LcQWtQjOXG6Oc0LUEN2WAC+l1IU9PnxuqWJR87ky9vy3dFXN0daKAOxv4Qqaia2dmD45gFew+afS
vCg0pHAPc225bRVBa8JsaA/R5hMeTVsU4tYUnnzrkACoewGeF8t45jR+cpxrf2WKQ+AOrbpqTbFn
uWdTfC336Z1JPzbw1DzSN+rbZlcgzCxyRs7IXo8lbil7Opv115cEdt7gkp6fuR8lFw54ApPPUF30
zpLR3bLTdCBHmkdzRvsKT3ABVHPAYSfgcLb+LHzSmhtBBstfJQBBMupzoLyA04NCC0RRywE1Zrgc
EPsH+I/6NEXmCLn78xrxWsJwVju+pDvpNSqBVR4df63bDn7goAOUNGKgGaHMrqC7GK0MgHPgnbjV
wqFHAECxcfO2IgSswIqbnTTPtOjbMQ8d1cXR6jSP7FAr6VosgxHt85O3qJH+cRWy1NJHjCNqAv7b
MePe6BnFQnSqkcdIQKR0GwyPQ2lD3mHRED/aEEiYvZcsqdOSNCsrvVE9tA4F+SWtRlps8LjIB+XP
W3Uuv0XR49ZXnBmDSvj6GoZ+mxDXMuUbZfrwMz1gUHtoyLSLdc4D2rJkQ7eZs40xKVGeINvZEH6G
9a33TpRNTN3M+Z2MI7g/aoPlY1sTPW0vuS+9y4CKxG3zZkBgNNUVH8hI75LmmhXhab+Z0PECITfq
Pc9zhpn1E/V4pbgu8tEvBVNks5FXPQF5Kmg3tzPPFKNIKBkHUTCIZOOyxtZ8BTmvwapFhP59JxGh
WfELbns0SUZA6BQcunLdyEWLhZkuBEkKihPx9moxqRTf8+3hzo/m0gnEmljgiJSi5e73Fj+HzDSk
gWugomjIURqwX2VKnXufwfhFOnmPxpnu+rDCpc/X92xEmmIX+PqJjEUyCbPPO8wgaa8SwvsV3yxP
d8/qTa/KvIaz4Uklac87YnOi7BUEfI1NEA/eaIGiP3ARskUT3rIfgo8fhRhqArQKeo1t1cy/vVkJ
sW2Wtje6o+dQZVua9n5Ky2ozwLBsprBZNNmEGiznCCQnv5Sw1q55kSo5ocfxzcfE53BtpxkIiFFA
JLioqVgE1h1LhQ/3Cccp3OliYK4DEyrDBToXpS9LNcxYPPHYhf1Bje7+n4HQxZgi2eF7U3fGaC4P
de3otpGW3x8ZyGVkJZb0aDNQnPdzR5LczGgfUnXKt/c9b0zt32YSqs7PgxXj8jzo4yGTOmnsBkow
WuTLaaEKSnN6ad6yfRAsdl6irGcvDFMDhfNR7VWTJy6Gtntu9O9eu2QkCrGV3yz1CojikabgJtII
pUrMnMSNeCKAP9ocFZqBGENHXf/whWKYlBJD0hEiEHw6jrzLIhNZuGmcR1c+sJqQ4gxlX252NTJO
x5125ziP8Iz3O/5ec+Hz+WH2Ec2PjksPdiGUaM/5W8csCyTAebiEB/ptRmVquGNp7CrwWXKL/tt0
biwxDJJyuMDfWp578l9G3HI6GeyUNcU5rU/oBa4J7Jc5dd43S547LZHnNxXYXVjj70J2Qrntye0n
k32yYna9dXtLcl3MkxMUMKCB3Y7lbPPlpKkP6BghUTQmqAxlgsShG2w2ZARv+ImBzQF/0c8BCAwM
5voanb9lP6v3sp4GEoKrK4uS3n611Gk9pd02vPZxlw8Xt2UVOIycoJcOIHYPw+uO17le+hJ4MdKh
v1ZB3D5J8n5ftSUIF9f15K+OMNpW/QiXLf0ryYu0KoPR4mj3ij+1NmDT105Aod4Hjxts9AYJROyO
xkcSS2AMN5Iu/FQ7o8iurgB4pE9lsUDApPnaLrXG500NTDmYTOMmkn0HtYbVOhgmxJbSrVRL6wTr
4t0bikPh8rF+e4J8dkofuuAGyCgYAC0/3sBQB4vjrScYYB+q1gZ6xP4Gf3vpBD3R4p8FOiHipqX6
DvcWJ9Kx0+NHawDMvyXvCV37VZqgpvcrtIPUsXwZycnUpa77R3O652VIUZoxO4w6rYtwSGRMqacW
Y90NfOg1qbvV4mOXheIwAK56N402UDWdqc/CyXiA5ZIpHSAFeM6YG3a4ldgzkmzgBeRgzGl3DBTy
a8iwV051DEQsxRTAymw7w5gAPN32MEdnY3NAMy84w3+KRBMuaoj4j+YDnU+3pm0Piulvd7SJEcwO
08jsB4j+FjpUvzYFapodH9QIDDHlD3JU9MAMP5iLTJBJgq+WF077BxvZaV35WTyc3qKbHN93GLmB
LDI2wE1MEPlqe3TqCfbo5ZmJ/St8rkQffZLywngo3h2bequns6CNWUPOl28VPyP+aKz++5zsEpH5
TO34mtoxDIwbfKWKiW5Kdv4lwQ4G8fvXghaBnU2nojZTYs2qR3RpvILCZ1YVfFc/lc7yCiK/2Etm
CtrBPOZJ+YDBYrhFuO7iJe7WVG2qsuZ6n1PIm+mNLFvNg+WrfXlBsZLHh0VuQkz+JULTgGr92Jt+
NdDZgQ3hwFDdITc9vr3/4CEytA61Diht1TU5i16vp6nvBAUChNfkxQ93l5TZyjOe9Q9FRV8Aeb8O
v+BBmx7tuqB2P55cVb9Dt71fzZt6cIPsZiYTwFuGw1Pw+PRVjlZbxCozykqA3GWY7TivOzqVPgv1
dXaCy+NP/3PRtphPz2QtTz8zh/jEajCoEyLUEykqDA2pRKDvDaoU+1vMqaoJZM2ybPlofGxTCrOl
Fz6v28rHdlMMquNvUYVumNeSTj6BU5zCs+cxZLRvngcQ0Eu/w4aouKzwcBA9iLY/nJuz4UjZroCr
6yTLMx35Z5XKf070DhF7x9T+spI7/pw3S3eoXqic2ESTfSYaUkxaU/Dkf2OX4B1nEGoYFOCIaSFv
ncNujhLKFNkVyZNZMw6FzfZoJMKVXlvkbCDcr/1kzj9cObPZ7z9eQ39qyeBupltHctRRGpMTHcLw
KpMs9FjRDHrBIxYUFDZ/VFOYhM3Ioz6S94E6RbPraxSvvW0EgovaQl/QpQp7EvVJxtoeNtFkUI5x
uDPKGZMhjfRtsYUPAzo34yGDd4kczwfX5AyuoYZkeWiZ1hVUpgfcyfh67NPbXvIA0h3hyPaYrTj8
VztFBjZoBd0hV7pN2HUMq3j3E7EKfYi25IcHUOITPdf9SwTwSSmI61GL1AkDxVO42m6P2SGM/SzG
B4KWm9oclvqH7QHVCMWkT5bt6hUpyYrSmNOzPjEDKjPQ472KMM6S1Ui0UxV7KLYP47jcNmk3hqjJ
nyMUU2A5cMUacq3J20c+sIKyMJYH3H80YrIQZMTNem3o4uJ3eW/sAefodT5gNMqHnBuM4y9/nZks
TlXGWzA1Y/wVm0wb5VecCNYtPUXjCY9uARbvi/tELXw1VjT9uwsTRJrvmXVQZSIwRmoiPvpKDzl9
O1VWQruGhxcHI0BJNqrzPKiQvUXUGbUstk24S/pUPETa5GlzedIq1f8LdkG3l1ifUgy+0zP/AqHm
qf4m/pXuG9O3UaxcgykJCa1EB5YrZArAjvNNopm0pJe0UiY+7GV3FCtIQdMApQUQAoXakppEwkGD
Y3VJXdxQ58+PWWyBOE35MMDAM4/hv4WnpDt1tf0s0vNjAN+6SEeAJlgDSiFMbvp9B1mhiYLzFcZS
rNHtRGH/xuMoc5P0gYPtJSkEKbwQRGPt18T5sMQHIniS/BrH97//CbJxKv9Zw/CkhOIlHe3SLFC2
HEaHhOxewKDcy5AOlWfuAGNz4MMgEt6U6PWUu7GC/CzKz6BxSNOb+XZ/MlOZjP6eQz30HXSjJPhN
K8Mi5eArzqNoaqbCs+ah6qvIwS7KydzFT2kii3vo4Zt5rvwNZjvNRsb2R7ivuDozZQf0KlRZEKai
WkOItHaUJE4PjdbKu0nL7DoNWugqVxGpZMm0E7OGNciySCrdpfZ6m6Ms0gQhkqoxOTBXE7HL3JN6
3UcDZggiSfHO7k8y28ylpswwLf3FFyeLB4aDpLzsPbt1VRNFTN2afRjl8Lw9yuNepWyrAFbC2I9J
I2u+HsfLZKEiBFAjP5XhFo2Ag0znhDsUc1zPZEjJ1Wq458pzzinXXe39kPA5s/YtM72Hmgc15ll/
ywrVknKtkx19yips5Jm23mFAjuqe/ocghEi/nN6ovtog1V0bGOyuAb/YS/+jExu2zHk46vWvn+is
kTgkajMF4UBKmRzkKxopz2d0BUYd9/KZfEUIaBFJ7qLCYbNVct2zgmw5o8TjKgdQXjJJ06adFIIC
xBaRnFSAFTY4Vp/3ism8qc5YdFPm6jJGC5II6fkdbO2hSqY9Z3r25O2sRQS4yJ6qX3G9g3jgC9BO
re+rXp7z3tM5YIZTHeeGqF2unNQpaJVn34ZaKf0sJQshUbaTxSRUXknDxKtmq60Ho2QRevFEG7Bj
J4Vph3+kq84ry7C64Nuk4jpzUMYD7Mhk+XuMPMPvZU89R5vPJ41V/Ir7LrNCkWakIKsJXzEyi117
GBtnfsN+1EIyNRsf9UR9Rxufycq7NOZUrPatBRWYy8nAgdMkKix4ubqILPfV//o5LzaeYoFTMZTL
s3VxrhjUQBDTGOrAS+7tRsLTztZefSzJU8DDMqTUCmBk7uA7e90QY8XPY/e8J1nIfe7IpoQfC5Gt
b/OozE1P89fjOwWUmo1WG2P6/5n42a6gLg8OK6fxcOy4xvi1UXRC492nB2soezncHblXgGpJpmUv
8gR3K4mA83MOJuL7iHLCBpXLLZgVMHwrS28g8nSHm8lQdXrvH4+7b458GXdMImCi2o519lwk5As0
OKhcWIRwU/mvWt8IK8CaotyzZ4QLzvZSjYP36P2ntWPXn8vhD/NCdY6TsCYRhoTPw75TL83mBJ1m
lhVevNez5LUTGNXEIr97mXLyVkYT304SoeEDN9FBed9VQ8bDsrEWxd93kZo3W8sCf0yoK+Xmpi8S
5gjTUMSGlxRXQKUvb8AJDrtwGGQ+wVVz+zTs926ESxtF0+ac1DxD0CS/EjS+EgaEM0SDFETUHH3S
msgqN+SNMqqw4x5i2GqLE/DWUqrA+e7yDxg+F7uUR89QQwr0h5L2POUqLuptFe4yVkm9qgRYIUif
rvG+b0EF61M7OZXrILME2UJpg2WTTMc69/w4hzBIyZwuZZsHPpsFhQSLiUebj/oRH7+Ey91rVRUy
CVGfJjvBjiEq1qt3MsJ2gTGxY39UBoi2QXWRmgBSvybdlV0uiIXxdg+wySk8IU7B4zBRr0O3fbUg
E/J7zBkXwvGdUmhdbNCD2DCGElCpsdvdWrJfPAeH+eeL183edj71xoUjziy39gp8Iv7l8d+rJfxs
1mdKAOmx/YT95ZMkKYwskoZ9TpxVT1GnWG0wy04DU2R3BBUYIwrxTsZbnk5nIco0o8KyyokGYROx
yJSrrBXWqcT/IAYYlu9PXviqtyMY4NhX3tTlabkzFRwjsRwDbflY4z0sOBqKJ4C24D9esQ3lPAbx
c1COvQvKJM6FZb5Oe/xApeadaZv19WHzS6D+qDD7Wo7mldzbqKZtk4XdTzP71DlNcAEKhLDyisGp
uQ7ZWXYarz4wrod2xOOchVMxvXZKfLV19GiswLTiSSQtATEBPcGZq/Dxn1ejsVdlUth2IaIZFsmU
R2nQxUpVcH52Mbwy0/jrKfnl1K78soa06lhnLvOoEVPRCTACm44BxE9jipirMu/C1iZoRNdWMdK+
O3G6j9Xdl0gIvo9S6eAPTGAw53AwqcSCsUHakdX5LNK4RjghV+NSqNbSO5IgiyEgpqbRud2DlvdB
j9lFoDMeBKIx/jO9cW/0+wWp8BMmW3LROXgNpLj+QVsPxaTK/7LzmAEX6556PA7USsxJxLPjji5r
OGCMp2apc2629LF0xadQU4btmWzU9L3DNR4J7wBHAZix26sdyIHUYONB4MGBMCXwwxdtgL8Nx+NB
OBqFl9ZwApZ3PF0lyWttau2bZpEBDpxMijFduA+V1WlCS1GmDhBOTVZTNBl8wh8b+F3JA6PEH7Ah
ED7Cu6A1hXhtghJzAnwoH+2+yRGPqJk14UR1/+H5LMpNVHdCZD1TZ7Ka2r6YcuacTlfYVEobd+mz
CFv2UIll8lCJ1wkYSMo8nIa1gSGn+nsLvSguOe+1JsASSEdV42ELiynOIAxW72AKcKLeU/FUAUg3
T8Q+sROlqVt+FY7e5uQA9EbHCF/d47wjRXDNfXfj5bTqQyTP2r/p/q8dNXAjLSk2lHNheXzQZV1a
mGJduAsIWSpjPRopr/KpYSPt1/GtPWUj8CWkG2z7WapxsskQ7P5nbEfmfnEzuPp4zdogjF8H8BeW
HP2yhtHHPEbzA4xUwtifHkLlnWgGrdq8l1Y+0He7gwmoSZ/9S2MUVwe5FCPjvGVcqHblEHm5O+NL
YEB8KpAUtqMvb0EjCmn62EYAhGdhYz1CjW16yDFlHYjGP0rt5byHymzxaJv/IODwlRh2NAZxVA0r
3a2+BYz3hu30jmBZaGlg9nqWYmG7vmMqZ5LZSzFGfGSunIlrlxOQYG7xgKWw4lS3K3Wv5b/8EUNz
mnxFxzFmERx2JQMeMcY3e0CGP+KvJyhDWd0JMr0eHRmaMnICfiRrpfNbRidoRIiATh1lNwzjzsJu
1qtS12VgL7XNqQVgb5xutSukYaASLCX3ClEE61g2ktRbGPVR2Cw3pIz0R+nDdew9wE99VrMoL4Ec
wEbtTCzA20mZIWHADC8fwhyRcJGU43Pktq3xBqKodb77Qx6t8Zjkv7Z0gMK41qjPA7QiUFQ3DsdP
aUEFGboB846NVzm5ejxVlwJ9sdrxLEPViEyyei5jmrIjBbZhNqlwwS4mRpgDdnjvnr9X/lMpXqmO
70bVFTLAewJetd9e9Syjg0OBZg5aPkupQA3AO3wfNra4cVVURHYm9uTyrunxWCK12s1n33RQCvHg
xQtW5l4Atz2ljlLYn5xpy5wXWEeMjBZSTPFGJdWNjKngyKY9/Hy2qEr3OwmAkZ8pf1ziWyozl+tH
aL2L/SF8UgpdRb/QyhMSv7UuHhurJsk42HQD9bF6HK5GjjFl3Q6YDO8Qf4OLG57jifqKBaFE2TBB
qU97/VBBWjPHZ9R2kY9Qpr13sU9hgnSytBBPLIaoE3UITGqOpextg6n4v7eDjeRvtYIVel+uAbB9
6WCKIYb1qXY4+tXHZxP/CyXFq9bqbAKwFVOYHMaLX+W3uDb/D/kAHkZwnOstugVRHlCjJpgAgm3S
dEy8mZOaDTGjAmnte8e9U6ubV/diiU1u2t4bKVNrIYsINHspocMe4hghsdZhz6Dy8djdQ1Cra5wI
UP51KUM81lzZgDNn9cARInNzjYXJRJcpJUg5UXn1iYaEykp0qwGLsjLMmT3Inx15n1l/koG7ddRn
V0G7IErB7L4JZhGksH67++p7ItKm52hAVK1fp0bxYEluQX2jUvIn665ljdPLL8U1r3+ImKO9HFpI
U56fVE4IKLdMiSFfzV0FN7tZbakmmrbAu+njXjq9SXHlK8mAov+g0wyyZvhThW5BsJ8rqg+RrmbX
fiUbxW1928ti294t+qbFZoaXj54yad9KyH3I1TPgpN7v47/9YkETIZbWMlO+Onuwd5FNMqw/Ju+n
ZKRG56JaCBesU02ArbudiQTxR0Uz7GrdQQsgewPcQaZz3wOA3VDUbAM0E0v20esNt5d9xxDdT3PC
V2rwvJjeqv5qX94IPhI3W9LoDDlzqvtayMSLRlp/RBqlXGKsu2+slqQSAyMweTGz0RurU0jDTAgG
irGgIX/Mr6sh0OjFtNqqhdjxyDenZF8Ol4YsIIyLX8FE6cOs3iLQ7UDFXBc8JjLZHOpWrvbO1yqc
BIjA6PvPaUiMugq7itP6V1H4EqttMW3ZAHVjPlmToZbjX2FacQnhU0qXwCwpotjXs7xn6LSJABq+
qX06loM64aKOx+hHozfBGLoFzj7Ioz5PyDyfIU+wHmoBHjtlzpTiuSGhvn3Sy+Kad1PB8mPTEFF3
1VXhcB8t0IsN8eLb54pMDT5c8UK5k1W8Ir9mFLy7cwZedCKqbRALrHyRQTXk9ZI0ePJYJAmErwGr
xV89WyX5V7iT6I66pJe3pR3MALobkc/a02JzJ+4f2YfyfD5u9UFomRDD+l+j75UQrRXNpDXDT6UH
zrv3RRzVCw0VmoLCnSdj27lwD335CngKTh29bOBWwxzPaftOfWp08DqkypjjEZxMw5zceNFIHDjG
w3NNRLVl0m1F48Hkt46zd5rW0Z5THh/YmvrGD1RK51penWuZGW1mB8fXCuDqb1yDnbZe5R+FLbKS
l10AexDZWUTefw6wFC7N2QAp8Zli0tDBiqy7eE2n/RJP1jvqG+VcEGBY3yZxTL9DjDUmRl3M8Uv+
+sxejm5z3MqtaP1WOCr+AVfSnFZLZ1G+d4qi+m33pDoY9eMOHpd/ggcsLRJswMFzTG1VVaE8qsoo
XEC5fdSPPTFSbCSl2eZO3MunxCIbki9sIbKxUzkZdfsdKORWuJmddwxGY3jPkKfdeYCFF6kseKVc
62npG63dAFo4k92x/ZH06x0wzmvcS+XUyu3Lki1bEpmxKtY8syaKovDnAA+DSpIGeaujfxRJVo8F
uTOgCnr4V2odWClKhDNqqROFpPjDgBRW5lmBqEV+yKtN9gKxLGHJo9vmtxdbdPu6O6lu6zQbVqxI
MEKIOGJUAMQFz53x8HP5naNOdFKExKsTcWfOZrLfGffMaQaHC9S9eqsacZSLVUNjCq2hnxmNtN/n
B7xQknN+jxEgT9UuGyZVrQCmPWDJyhCNeK4NKRw/1Fz4EVrkjhtLKQsOQnTmwC+zEv8WUL0pZzs7
ycw2HtTLop+IuDkz7mIiCNish6OgiJFGIbg8owBo+k8lw6tC3eH6gC4chba9BAI8s+EpTl8lKUuL
Oh3nPZlOjC1v0LY0UYe1GC5PgWAcqFhmV02se4Ph1ZsLTnLep7Hcddqv7hAW1JRsL+KmZao05Ogz
tJ3HERrpEIXhn/ndfTIYLb+ZqIq14DMEJUUMTO5YyaFByOiJthMtYdMpSI+jcJ+nAzXPN2SBQLKm
uKuZUJEwfoModnQ7FRx6sp4Kr+cVkn3vq/g2mbySsuf5EuFsd7dNm2c4I/p1XZ4tnm4W7PLOTNAV
jSbS1TtsVQcvKRn43coPl46h+yeefZLmgYu2MsLCoY+JftfGm7qyIrapg//42wTLPR8BV147+DwM
o6LNGgVJV7oxqaTtci12/iYeVomy69DQKRleWBUnWga28jQ3tzwHYDIdCPLDxT5HY+RGRHSQeRaJ
8bdEDdylZEdt8516/GzW7JArmC6z8nluYGhdXxMEjms6WSgRXEUmarM1zfEUQcBz/k0HKFhsPdkd
1nA4syGTF+YHD4MN64OwxOnomZmJt9qwXrFiS9bir6hcH7lqSLIQV5PlEwwRRjWuAaFp3M5VZY7h
OkbzXeg3boeww/dAa9yxmLRDagLjnNZHc72m4H3AJmoI0xW0JD34TEldLooYebJ1yLNMNTlRRtzE
L2H/IxNW9Hf+hhLjGZPo0SJXjaRmqTobPlpMtjv0r8vcE3K0ew2AkDWkSI/3GwbDVRkFopTnaSeB
C/qrUCxrkw21FNkeVb44QWSGKhj1nxtMhIe2VHDpoq8wr88PbAyccpocil0ZqjKijo9ikZHwN4M3
E90UI3HhcnPJcwZu66loFwGiJG72tLPQed8ntpdM5985w67Fs8vK/YhWoyZPaDh1Yle3Fo6e4TZ1
7CVV2lnArGuhluh7GqZbfRO0Mqerk66hA95doeqieRRp+QDV2rkWgjbD8zxVjGnuNr/1RWWRMgGe
JFos/OhT5Up9xtBQuHy2BTjSCmk/MzUoB4rEnVbIY0c7KNUZUWt+CHAuiVsaBSHawN4ow02Sr9L7
4xbVc3rqyLZBFvJdAkHobW9q+ny+xS5ruqipLEqjaoBLcAt+MAoZzIrvqYjS5DGWg7c6Kb0alvmL
5WCEOKk5/QepLrBOI1gx0bXsPVn+PFrjQsCsZbKMFaR8SNW30+CxnW2WpZ3Crq3JG8FDNgv2n7AU
m2iIyY8b3HPp6Wfcmz7Ds0QkaK6pnDYqyVQTVM3a4HYYW7kx6cqFGVruKCwtuoktxiC0f9hT/CME
dQWdeX/ZFFVEGp+zMpCN04aDFWw/DcwEwat7O563qwuvBYiMbF7dPVKPikJHRJMWna5v67FYHNYU
PwXoUh4DnirFoLT9bNvPG/VM7reETTTINzS4v9rohcfJxuALs6O0KhxZklYrrPxssvPtYHvFsIq8
Wk3EnKgi60H1iBWQmoC/lZNqPc3RDJPyY2lBjlqQJyNBNpBugIEB1f//r/87KAeDa+YOTcleDuHU
wJdrnIB2OnRmkhetMPMrrZFrU20M4G9TOZ24Q6Njzlc294thLkHss+9rZVzd0M4KiN0Sq7qlHSss
dBO1Y5o2bNlC+Svq1uUcWKOGpzONUoJbkrA0TA2/gaWlEEa5UaywGzVVipvDnXkcjHH3Kbhp8s8a
fAto9Uwf3wWSb3MusyutlFbQrhPTRobGaZBr70MduRyVxBY7bKGnUpipFY09bQ/oZ93w2keQ+7KD
dD5EZBa26IP+grHbm5fUWZHrTZLXzOfZyPPue/R5R91wm8oNYILXL1bXxPmRI9vbzcgf96+GvniR
X4Zo0EHitLvQCksHtzmI4Pz3L4tIj/6/W9d4lP5HNHFEQ/ysxC7maw5Bi4ID11fMtgy/wKEXIzq4
BgsqfkLSqatJ4F+C92ZrTSaqa1sc/ZmjSYnrmnmmwHyq6L4H/tEG+aNXKbY8Do/e3wbbKL3Haumu
Pl80neLgS8yvpINT8i4ylATAk8aB5eyQg3EobB9c9yqLT8Yp664233TyTfe+lNbf52x5P7XTXIUl
WDRPn3xFFTtm/eCqPK2hVQveJ/p1y0SRIqhXj04hN1P8isyMcm5LCAYQhXS97bzFxEm3Jh5m6mqw
uKQ7aQLJMAA+trhra8xk/vvGG4Zy8q8zjjR4X6cehm7uCLak7Ru2v7bD9+pNrtLR2E3/8Ep/rQKe
uG+l2vujG+llZrQrA15RWpkUQdl36C5TWRGX9kqhiUaU8tR+Qc4C+KPVf+JRpC3fS6Z7YwkhsSBK
+HD4HClWRhibksAzEHl4qzG/isfJg30K/pUuWF0q/SBNrgSXrAEZf5nFYYCoHe5HObsRQ7slEU0o
574U/pJrd181iTSP0YVwccSJa2tkL/oGiGK3i5BH0Qr1HUJfjxvbgdlKJ4g4k+zHAbVNWFwLgD16
b1x0Cc6Tzq9QprrfLy3Dzkd/w8GtEVSrw4wm+a9ceZV/V5kXMqu7VraPM49OUqgXQpfC565hjfF9
IFP0v7mhUQSxXWi8O0W4a2QeMTyT1uily4tECtkV5PcdrswbCYUCNPvu+Vjb2JMyp0q4Oc2JSFYQ
YtSLgv7lZ01VicEA289ToepvX0QTKuwvW8CeNN4Od2i9iSlJzpbn7J4wQIJOlgEiRE0qfiJ8k4Sw
c65plkclud4H1If76F88vsJy1hFW3YqR8jpAhS1H86b7Vz3EU4W2OSCA+Otpxb8LEYSxUFWTgjIT
0zpKQSYRgZepO63lucy8IioSykexlER2ZkB+crXs7rlX3nrK0KMUm+wFW5znG0+mEs0cHpgKO9Yz
DnFyQDi5V66HoqPn34WiQNL/Bvc2b1dLpoEIsI2xNoFvkupFHsXyZGySI/uDLLUjBMUEqFd6d+u/
rMklDHIgqrY/EvPswj7aKeOHsSNm2Vzg98ZVLNBgpaQvwyHF0DpfqonZkrqyBqvZijtpqo/ILufd
qNCwkJ+xEt5NrMVwxu2OxpUJQEC7BBNbtM3UbnSHf6MYOs3zct5alvXufjMePMZNVQutXoFs8XXd
q0HrZAUx8M+wI0UsvT1hCpegcspl93GYuFyV/vHO186ZTJewjjrcZqyb27khMQ/B6ahb/RCgglLX
wrdDV7ZAeFNoDqf89AN1gS68CryYixGNN5KymYOMCIDbmNn3UFxrA98v+4qrp1fk5wPq5HmXH7jD
v3mi1HZTYuPTqFGxueEbAhp9fCYeNIFPvdgGZhsUor13MD/KK1AsxEEJy4d8rYTdRCZk05Y3xrjm
onHdLYwioC2kTLEcoTXNMPJfiXFP8JgBDILgwRBus+Yzi1ZgNZvBnWDtiA+Pd14QAO8V/vNc+K1l
fzqeSPuun9ri38nOJf2rt3eJUYYgjnmdN1K/TfW2b9YoUpkfKH7crSefnuOnIjbr0oR29WCRt4Tz
NLSSAy6YmEafmeK8uqach9Auzs8vpW1fDMqTUJKyIGokkBLRAIVKgfJdkn9Id15gW3pkAkNGAhAi
JFopIO8hbNHb9PI0am55G6jg3YexW7/l7y9JeFrosriRLUnAc6Wh9BVD1jE80C9oNUSKRRg367XG
wqH5R3LnKs8+h+pjW6qpjEVjogw9iHfvA55Vmg/p+dnXCLFKbdXQ4yqu8DLVmXU89hWddg9eh+PJ
2znnIq5yp82Y6FxFaMz0VZq1a5fIxQK9+7lc1LSk5e1dGf1r0xSuMHmBmbWbySeN4JpT1EBB2NE+
EtXhxgEn8OwOyPb3Tg6JA3sEgTZ3oAvhzX+wPaCegjZPritRCNbEwRNcZ4IW9uMmKayojv73SFy5
z1yrvCGG6wWI2QTnN3YoUdMIT2h7IXe/0CwQY0kgKeZx2jPLjnbwtDsHDDfNHlFQAzEUlVPZAqCJ
Q8Uc1+DlGeG+HGAZqwre34pdFcr8LxF76WfKWj1sYn1Tk/e6lVsv1ge66TgATuzUWCljv80TPEvZ
hMiH4+eG4nba39BjHD0oI/X9jzRFXVucdJZncMedJplTijap7Dr9MLnIDg3EwOIkbOQbTjQl3OzT
J79zImBaQebV7eEPMxhGJg44zKkngMtf+ynBFvUrk4PghmKHyAjL2uTWvM7f2M0pYTA1gHbhuaas
SonEiSqD8p4NuC8OxhLHDVlJEbM7H6sTwxOOAH95xYwtM/ViVomVI5BF8uN0FZci43bKfWzd6MXI
SBLSSgpPOrxwVSwi5XC8idrcC2wQ+IOm3evSdYft/d/imTGdLYqQk0GMSlBRJYG5uoOD7kEv4Ldo
QVmHrDc2qszO2+nAYzNCXRfNWfmBHsUyGrka79rbiL2y5Gl62oZ04CHUAKHfBcSK4DHDhgo5xS3y
q0lIRa0qkYwB+G4Fompen6o1osINJetnJjB2hL4jRVGN7HYaDReN6JYtNn5E8Np3JUu5qhZb/x+g
iF/MIXJE4eYRhp2pu5h18MkhGOd8WGbceqxL08lVyjCSPsPj9McAUFQugnkRf/WYaYYVwMLiPpmj
NiVK5h52r8Tl9cvASaVA7eHbZWD+tKBJoCY9mprBjssz4gToAL+kmPRNxZ8hIW6Fv+KNGtfj5hp8
qqbgi8mWVH4J/LhMfJOuQF82E2wdDSGgDqJeTlFJ2q1OPbBku7qk9gVrOWwnmzGCwye2kdWvjx1L
TVnwOzP3DjUEFb1M8XJNxEVJgg0rzvx4hKiudVb7DFEJ7QUXsEQcL/7uoB1R6FZ2L1L1uoyKZL2O
dXk2g0Z+Ku7XQzUecnECziJdLK+Bg85fTY7dI9AtdpC/07d5wKxtreUM28WMlidZ005P+3FRiE0I
ehxgyjKoU1wvSlctetPT57RZVizh5NvskZosJ7b3ZyIyRxS9vEtM+QNzB5KELVZXoOiCcaxiwdiQ
DnsG44KovqD3jJ9sxK9zVkwWvMD+cxJdA8GTycPsb9eqCTO/6QRMMJyL3NBu3TTIGM+2/aLD5l+a
zq1MPA2DMhkCujoONvwpsrJA46KqOr3DdnALNzs4+JMCmcDsGsSzHxtkc8fvhym4I5AZUbwYqoHh
Q+Bjq9hAiqUAqyfpKtvZufDIKzXQhMcHkdraAxEp2kwum8OYDeEHIQdHwOEEybHKmg1zf0uZRyP4
qhNhmNBqTmuHqCEXAGkhQ8hudAb0MhBJVz+4WW4ggdrRAnFpCXz0uGCFURJVdi7PE3yX5U2cuUEN
1GCyV8hQ7yhckDIgu1+uNHkhrFh9Do072+KOU8wK5nhM8beUkFC+cnWgi/SA93H2fIXj2Q6ptnl3
D5MXNvFTJgTBgKi57aunbFfJgH5F/JqWuRxwEq74V2TIk69HFROCv49fIkKuDKZOavmTG77q7Vgy
lbujh+vKH62vI71ZWZVzoOx7g8hBPAyMf/sjGHeJzS6ko6EL+lzWZ7Qghtx8aI6mta7RWUgyTcCW
IjUMzW+gS/+3zBesQ5FoJ7/74JoHSok/3w+HHaKeBTYmow/KZq1DEX4Rcv1DF9hD6E3mala0BKVN
J27n6xXANCDdCadG6ZHES2jiDBn/7peiB3HxWTKDstoqWHX8HvQl7659N49gKW400U5wT0rd3GjM
xcBrYUGIXkXQNE9nQgQW9CdNlnCgWFGXi/lKQgsYSBUtC8Hb4x2X2Sqec9fVWwQdUyuvV8ArIt92
n53I4UY5cddSpwcqAMdh6hZ0LJMeEJ1V6iYUiPbegqare+Xh2ct7UhmABLFlv73TbL1ceFhdbW7q
r5Sy/xZv6sN2y25LQbzfWwVY/ttJU5TmyRqDmgGdrGgNiLsFR7TGqg3tdzLa1RvKZkEzD+d3fY9R
eOazQR07Irq0TyTD1Sxk2XAFRoZZ0/XiiqL3AczIL/2q+lm8AgKMYV4GZJpRXoV26xKMU7Lxk27w
Bm5qRzRz1jjIyCZekTtTeynKW7xHQ4HYWWK/skjtsieWtuNh2KO4HNVQLywcwR/qmR9iL9zA8ON5
3IyWWB2QIEzE6e+t3g2s5Z4DVc4/HKHGNtQgBgZ8jYGh9BHlNRLFwE2dl+svKuodqCDUoI6eNMx9
Q2UXMcyckSkjPhs6WaQf9kdJX2NpTRBV3zh/4TG4kjTgQ6rmCEf0GjGiVeiDPLzz+fExMRPREF2F
15GjxgHNU9YJy5JCF6JhXSxxmdkjYkqSgiOzdRjwB39a/5IqO4KTAdFEBTKpl5XqWyRGvSrrDIWD
jD65fK/WYu90i/sbAf0a1nh85OmGQtnbaJToYH86gnyBg+tNsC0LRJmhDrYwBIr/7WAf1E81U9La
BsR7pQOo1GAc2kSnRsi0kSqY7UerU6ZV/RCiI5jkPZGJT8LjkBj+ghAryjyH3sBx+yy5iA44Xs3l
C63IAEH10O8+E7s3F2tTIf7EAShEY28BJlbUaqIbWLhhdN+ecP8aRDoOF+JQBq8T+z4elVbCIDQV
5hqqSK3/ldhQH8oymMrHza6pKyxONh2cZwRUORUhCxsWoTR+BrecccMJM0iC0rhDtDBCjbT+nnrf
zxMBy0iGmXpzI/6A9RVp0BoO7CGbk9a9VACri7eX0U5EmI6XmLvMpTj5X/rsUDWYJf2AK4eh2tcB
v+ll9ghTeeS9YCa+YppGVsZNCklexGkUAIQofkCVOwv3WJI8gRx5GneSTS/KRmcT3xcK63L8H07U
24//7ZtHIzKyiowtlSwf2lVu96yOEW4+bTa3edDRqr3gFRuAGfoDY5UWYKZTikjjlG2WF2HUArJ+
1uhWhl/j+RsyhhLQh39TLqjwYCbG2xMroF40MC6b3l9a8Po3xchjBO5+XMV0GSJyz5XiaWKnJWqU
XdASaU7WioeS7V3Xxvc8dVK3IdznBnbIDUauNNPr+5h/LI/P+p4SX8HdQ7OnahZrjztePc93bvO0
Xl8zy4S7N+30Dh2f9S05JYC1wv7b5p8m0KGlbvGKGh8Sn2pLahzUpMkslIni+vahEDJuTsFjX2Dg
htJQ+HK0ihzjbRL03UpGbECA6laxpHuT9XaIeP+TbL5eom7LVyrDiqtRm6vu7lzrR8ZIljM3kZim
EKOasqH8tfzK1h7UOqKWOwhDQJDtBC/ydH9+23UOG/Caeu16Nfj6LxcLr6GIxJecFI3IgUn2oTwk
MMmZ6eRXcWxP3kQoDGbr+QQOk2JXqfyWBQ/oVpZQOnoYXKx8FHmMj9+ZhM6Ib8mf6oJidLgzrLmw
bmtnwQnIr/sCg+EQ6uDxRwXDYqsxgd1rKkhpAJsXxIzdxOgbfp9Z88O8rd35LCZkUdYAgL9vp/w8
jOa54qLja0yXt/Ts1S/Y3OPJFk9o31UyXTbUa+b4oCV4mFyYRvs2hqb4BaMNOET96rJz/4MMRQt7
LQq6WfR1zX+g8OsEeOg3iPrNLf4ssyQlGoNNdaEykZmgXRo4q32jb2ZCswAj8kYJGL365Do6q0HD
KUHSP5l90QE0M4zJmsrQMVHWTyA48L4IEpTIfZDwyCqZfi3pGqUgAKqeEgwZeL5VVLmoif/630y5
RrmDezqEEO8SO7nKD7EnYVPx1jCVZ3e0gLUTcNBHRUOOVgmdquwLCPWjzrXjmbbVCdz1V5CpOfq0
X+MNudUoa4UZIsneLyN9xmdFL1ql0G1eQOtunoiNkfYZMzKDFBaerOSy43WZA5/KbkD86IldrVaA
6YUjoQ2mPjsiqVocNJFIPAMs8V3A8Lcq8mUk+sUqhxZty5UH6qCQSQ2qH14WL5wBBkTbUj/cFNSP
oz9QCK7urs6G7kcQpMisXzkbZFzv2SdyF7p6TfJ0C5Krv4yqt0ayz6EuuvdFUpqRbcju7T51iuVz
SUwT2U22X/eAST4dxVJitfZ2a8yZyxSvAEYLVV+LPS+krlyXG/7IbuPziMkC/KPfosdmJgC2kDlv
4SE06yEsSxYcwG/6JfQKXOc1uvLD68BBKDF0qlRAsFdqLGf0X9gUBo+4o+fV4aRYFc0yA+142dKq
4pyQmPHBoQISDkcEX9jSSm7XEDXvYHSQNvjbzQQScAq5AAfSEwArRgF2SIKCuN1tMyLxeiFM7gGv
y+nw0yx7RN0hEHX0CH/xDIStJCRQfGViuOg3zIc4dioRe7k3CvW9pmxtkNqF7mEJ9paZeBovrH7o
zW/ltmevVmg8tBuFZrwaZ2pDkCQopSbXDoDyjF3w7kkjusUpDCh4GByKKXrv5CI/XryRgSeuY8iU
X/CzQNjB6TRLSFClGhRuBtZ1hxCvAoXsMNuB3wMhBev9GC14onoKgRJPDz2TzxOwKmNtwIcJ6eEf
8b/n8QkjvG7V35f2LvkwQykGiRmjL2leCqqBfrsmJ3IVJFZv3R+h1bm39mT99PpZiJr5oGh6QVVH
CHJ/kw0ccjOM1z3vLEz1Fdt6Glj7KloV5YBDLFwG7xexC5CaK53Va8itFhTOnqNGg7wg9XcrASxE
Pv0krQ9JEyqch2lLDDLyVO3SQ3gWAtKt8Sl6I2JdUDcBAly/XlNOpoGA8l5CJs9Fq7v1AFLjzsqH
YIjG/QJ0eE/wI1cwQU8uOLcUUbFq1h2BVjoJDu1KhkX+PsZ/mZWstRliEv5+KbHsRxhQVZ3HGc1j
W6n3pL37UoC3If1DnI/UCda3z1JjrCXw8Y7QZnfeso4HLrnMpY4m4jRc1vv1CME6Dx1PISC0yF0+
hF9k7ydtu691w1Q4VWazTNWFog2baHciXLilnSYxbbXFaluo3TgHsDKxrhUG2RzHwc2OAXnGqMLN
BbMm9ybgNWsnejM/sYwgEaX252IN7gLU8ah9HZ9ZrwcpFiOGZFGxfS++Ol8ZacMk4eco75yJ0fXL
39nHg7bplzl+qYNWJDpGnQTlRwPk9dpohA5k42c5MKC7r72HZM+VMoYWYKyBIo2DVzX0SuXjaZGd
uBScB0YRRKmAvA1QDA58SBm+K/2ZDAQmjjFCHU108qL2OWkG9WAb5zXVy5E6vYr1NgTwKAHFjFNN
Tafox6P2fU3T8qrHTSxgdmaz3paPoNZj3uUBBXX2drDptuO0IfW1Dp3/iz7DVi/lGFbEghteH5a6
h9OKREVoZf3dvyOub8JJDDj8kCiLRyZP2d/qjQun32it/uTwSE2PHcZ3mACqFZ22LR17PXdKzy71
1HCHG73fHubM829J/MnId6AlbZbMYa7y1OWm04xhuSMO4wB3bRmhz9ASLj1YndYSHJDhfUT3eIxr
Fx/8FtlBO9Dy/WT8wzO9Mr8e5nE5R0ebnKKXip1Cd4qJIEYgr5JWsJsRaBPl509XSlPetG3QvHIj
plRtOSY/rqwWFi2x4JgIDOYETTxLU9U/aGYmKbxllxg9+67nNzfsmpuVrKlP3do84a0Fr4SR7S8/
XnHHAgA+pLgBoVg2Qq7CMkRuCvNK6S2Y9UWrA/wS5P66Y2kl9tfQ+o1xf3/yzC0NuS4K9ztMarYA
uKg+WFnJb3pVbchNZyB11XJYSeNBAsXHEo+/Wett8AnUwumxOeCBe0fYYj419UfIcRqWUobVqeDJ
4Vv6gfn+3D+I7UdUCIsgenJE3NUE3vCAmikYdY3IzqiPusVtCrJlzrxeOdvbT6cTm1v+u4ml+jNS
j8vraD+op8i3YpI3RdWQeWeAFnPR01pDrcTJhjHocb/k9iCJLF8sGtbxOyKKHdmP9M2dDVfPIWIC
q2YPjQH5cHTeM55vMIU8KaoUw1O8Fli5Lec9aoPEc1tp6wjdBKPDznS1/OBcejUKWR/sajIQXm3f
qe9XhaA6MR6rwkYhi1+eUJktOknjhpbZ4WxyUGxJSbg4hxslHAQ/LxPLMVcCvCgORbqJ993TsiKp
WJVx1z1Dn+XSu2y5uLPi2WOVKPRCj/OvRj1SNK30h7kzuqAkj37AZH4DvrQ7oHpfpqnWXJqI+v3V
4LKo55glDRH8SSzmD0Z82bz2khOJQ+FqwAPIJzJ2c8x5SAz8y//6pI2sgrcDD/xTL0ZvHotps7+t
JBrSl7j2PqXWjVupKlj54AfVxnuXOzl6YlSmHzXBU9Nj5gMusJU/H58BfmyWUIucPLnbaG0am7RC
6JlO4+7ORXrKksZNLxEYN7sT2lqqfLwz1PBqxnnOUQHgg1//XI4IEUQnBqFhsbBsYNF+MJT9n8xv
4Phd0dSsyFIySlhFLoZEqFvUUKZPS9p3arxhuGJOvvrSGUNj9GvVRzzYRhC4jllanK3BzFx46tal
+8919PdtA9UPMMyoFDDdgPJPnLa8UREP+Cm5lSOEFzhM9MkU8RkuKU5DbR7c2OT+bSs5ScUEM/7B
wdx8qN8GdKwqrw9lx5vP/uDjtYwDlOCoTJ5uqqx/p64/f27Yygcr4qMI0Z1Q7Y4+6wBxu8XjF7p9
bioBbaQG0KRUdh6SGXE9WEFUuxjbCXqZzWgBl0jY/o/Ds7C1Iv+/itTqjPRUx5DJ6VEdoOJxBp4A
B+IARiwj4nfSgjIX+j6wDwA6Ho9uvY+xLDaGiNU4xotvpoUhAlbs0ZPghoeUFwaRBWiEVGj++eWb
SzmVmRo2uwovHjcP180YF0LRv5knqvEXI3gPnKrUOmRzrcDiBUz94oMsWgCBMMLgWc6IObZov5pV
HL2NX6lrkAKpSDpD/mJeam38br4s5uDQcfPn42s3nq5l+umfxDzf3B5HH+k05SQn/kiCF1oVvMX6
iJY958PAea0cDlHT6BTWHX2SLrVuEpzzaw+o1HazHE5PlwTlsFwhuTsDu3ogIdh2ZugDrRmh78p5
PTtyciZFTpoMd2HelYn/gSDSMcO/ZqjP0kdgFE6MgANYQTm1JCU8OpOjnmj//t2UiEB5QfLMOVT9
q8OXccW8tLod1uz9/ThlNsorsPlhfKd+3lojzF9HCBiTVKAlbtUgjY2MJZEoQYrvkoXHx2GArJb0
bmOxQbXuKXZFTowkPrEqrk8Qhv0YxghE51TZv99gjV2NG+OyKyV1lzNygsHgvgfvZH2Y3spkX76W
z0BFu5eJP9Lqa3/lNkCNrEBJQlYsCffTdSlh/x4F4uFBK87P8dhlhgz/9+t90wLt/6zYf+VpDNJR
vzBcAso3nlaTsGm7FTxCNXihmmCMyoJxZYB5Y4R/5b60pQQQyUgjZbZPdDTxZ9NLBvWNQbNcdeSl
kEJqd9GSaoUZRnGBNp6Xxu00kG3BaOfenhUbMkhFAUPRFOw1WjX0oHZGjGSRzkr3I75WGES0o3Uz
dgoZSxOoPSiEpt4H0iWOldkXdWoo9VAp/d/eaPltnw8AU+4iJ7wHxswEJ0fWv9nCDRi+oS5He+PR
Tajni1K8t3ZFvJPhzJoRYQb5C8rCaG0Ydm5qam4SFbUU0fFMS3qCEVPmeS9MgEUQDUTSgbBW5ujk
p74ZDQ2PRpmp7F5RvCi1Se1pqsHs55DuwsDBuqfHL7oU9iwN7g/UYUaiazfNSAvUxp9EU1RO8YbC
u5LC1iAE43VQSCG+pWurojbfUp6WPNbUVQcEKvoqYAOlbdE5IRBAiVXWkaFS1eOTBKS45qRzb37k
CUqvmkQVCWiB399HEXK2BwvfYYFUrxbjOI/ZG7ll3pDRmerjMCqf5bdJNnUw/rIci+JX3CiueqgF
6FxFrwmKAPwDOG21veqc/9xNpvOMBK7MhzTYqzjVkZ5gGrg36p9a+LZKeyieMx7CgY6ltjRaOaDv
uFcIUxbd3erlKcwI0t2IubZZknujG0OziNHdxs+4phukpjsrQnYFpEpkby8LBx84Rk2pi/36ARGT
RN4+7eINa/G15DNefe3vILPW540h7xdYfD13IWLVylKp7X29865wCXFwL+fyXu2m169mTX+2pjVp
UZAz/rVSFoBN2eVH53zFdYZZiwP1Y3cTcW/GZl+K6nwBB5aykNhunDl5eN1TYfCeS7L6HbKREsje
OP+x2TL3x+ib/90rWZlPD2gFGUsYEKRptVxBWr0zN73hD2YLiaUnUiZ4kDbF3qXs7dqD2NJQtwOf
trGLc31GgnnDWtmOGEd1GvN3HyLJRX87SCFNeMbjScIvtvR2RztYGLphdrn479IdYEq0tE+7Xssz
y/bw7/eHtZT1A0IY0vYa4PWjWJemrkBhh6URtg1uqk7GwSTQgI18CiHiNHKvg8TLpkqsjKHEhiq7
LVUfyBci0afDFhrlCyqXYHDwXf6B4SUG0FtS+WL+wyHmVLdxlkPWlvPCCwYSgFDr8icGB7DUri5n
KCUsVjq20KPCAfhWRGvNILQfsfzZoVE4j3OnbC9ZcoYEeTDR8QXAp8rc04WX0jr2akzE+18YlYhS
PD9/FloYrft7Ep4x2TI6vmfdo0OjL+KiX8TbpKfy+7QywiF2a0uptoYLzOpsvXDjZWpPRYS8PIZd
jyfjf8SSQdx871oElN7L0WbI9UW3A0c1IiFpRYG81rLdXusIYIOyMV7eOIXOr9XozZ2wwQ5r5ceX
1RMZHUFE8ogtnwjVNkDVCrRWffNJFtB46yO9FOAbJOWx3ZB7i/1wHEVnc2Ange9L8JqDkGXnhYCf
forpIXOG9p9YEedTBKhbCN/o42bKpfn508yCn6WH0Fd8ttiTtSEvMR2upzJFuzppoRH353Df8oxK
tK7gPSAER+kJPa1Aw+i0T+FcHa+c62AcQ50L8YmyuKVEBlIorQHK6KHibzvYPIYbv12rCZ9zYGqk
qplV1KbgsgOjV8vtb8gZb+RVZ7YByW8EC+Q+mrjaSA+AjN/hRGIyI1Z5d2xeH2zXxGGJ4/9bkfnj
rbol3MIdPQjJUyRYsupoqqMihdEEEY1NMRojoHACdw1SqoBKVOztM1vESVMdaxlQxQbUyFK5s8cD
hERr3Cc83qgNrXkm0QROqxJvYEYN93ZtDo6NYLA7MIFfXLIIQUN/WrViB4PaY47s6xumRVq4r/zd
Hj9udmy/1UjvtAuklKEcSEg2OpYLsbeqs38xZecq7UBCN3ENECrHQlG1cW+AiskYqR0trzT6uHAT
ROR497IUkUD/X5tq5VgsdoR2NxnRIy+n0Yaiq96+H5w7Msuski5HOt6WQRIuQB9e73rtI3CNY2Mu
piOrGdodGFzVIKYDyMC8acAHdM9KFbLzp48+FE0gwROJnF3xO58eAgiKgTk/5W9su1YH59Bgo90v
ecInrwXRkR13bye5p8TVSr0kEskvMOcDUhHm8gd1P3JCzEvzr0nbLAnGilk5jkYSA9dpUCAS4/QK
SVR40AwWNvcGn+ffcF5EeRkRS/fop9nrTBB7E0AmoTWzq2jrvnxryVh225+GtlxIw0eAUoRaSkwQ
coTI3gvdJHmIQ5dMJCiE6OlHLIG4Em0BIYVtr/KGpoxBlU6nLhmXEOotPpnyaaqz1Dm+Fovx3EF4
VE5vqDjqbuRNAjG7Bz4r6b6qZrxuqbpREpMg9UCtKz6j/VC0437YaoKg/CLVlbIIYYQ1cJ8Ng06u
n3W+5VpNGR/SFRWTczVzxM1URvVuVfGeGBgwUEKxa5Ubi8/oEtzA8uqVROX26ybHyfu4GTAue492
ne0/IuZhkeMp28Cxn71xyoK7CBMFHVPUloJKNDbhaXR0ux1NrYxlx8v9t5ysyhKCYl9wPWI3IDF0
VPgSSg91rDCwFpIFGiY2aOvpmwiq4/rqdnqVd8Nfnaaq4Z/gtIquMPhppkCqw/IzW5ixeuBl0yGs
7F0KMsDxU52iUrdkZHW3+677rL3fTGdh/27K9+LmdYOaH/lyW3Lf4yHLJ3sIzAVNO3yIfpBplcl6
RwWX18o80Z2P8Y/cFSqtaODVcLOrSJCfiEnxH/oI8IZ825p6tT/2qtdD4ypPDLvsPuY0Vwo8Dyja
dsRutNLqpCDVR2X7VJrKZFUI9s+oxez+tkbtyr5eLRG2XaIS/Wy7QHfni4VPzm7vqFCEDD/bc+j+
3H/CStvkmRYneSWeTjwrGF59kdi9ciy8a5+pVtytQ9YExAUXBLc3pzx7bSoDbgfAFOlRdqUEdjNo
MGFAANWIKFsUV2DjSxjI2Ig37nNCfa9HYAp5WpcN1ElDVrTdDLr0EqSaMH8JgIvOpoeUna4sejbX
LvSk+l7RFl9mV3eylYR4mKX9wRKOxxin5I6Rz6/BHPIop4faMI1eav/VsYNcKlEwZuS+3ytzl8Th
PUBQmq0GTXMLIH+JqfVz30nvx/BpX+ngxi2QfWiCUku0mL00V/X7ZAZGFKKiSouPqfpF1TwneIJX
Bqe1hJtaPgOl5ake6qS7X79QqSxMj70NiO3Hc0S6H5sQGTGdCepMG4HR+Y+h8mQXVW4dC3fdreuo
opGTN9FAS7a8IHtFQg6lJLoxhwuoI/YvSOBpX5R6LpCai6KwH26Zhi2jNorwlmYTJnH5WBKXPRhf
ltR+ZgFhmPYVEemJzdO3ZZiPCltbIUDJHhjqir53gdJbKLRkg6wjPYQQNfgqpaP/uSjBN4F2qiIo
XKP/XRq9XMcOiIKdjhvYq1iCG/29VDb7yiRY0ulC1mPSU06UTean0n2ZR8BrmyGIlEhcT8iZnFH3
slphONlXfPDJuJ/mYMuW81htP37KbQwepKHyKRi+0WwbhPGR+osfVNSBaODsWvVBEq1Ax0Y9R4RT
AyXOwX7fHfdWz6S6Zm+vIomu15vlbNvaHieaC+aBX3jMq94k85M+sovnOzV7WzQMXxhzO1Qd1yhs
YsmkJggQOmlGmV5pdujt8XbXNlE5Q1XAZI6EfFOnd49hFCNHuNt1s5dgRl9CG2uABGdC0UGpSoh1
/rtL0OYC8rNk0Ke7NV/d6R7NjNLd9IOli2N9Nqka2m/zeAu9A2eLdagkNHEtiSpwBjcte43wSppH
5vt/s9D3B6pfohAdHQ7AKCvaxcKW90TyURUTjUGT/1fWPLBpx4mAfSKVHqQEDC+euI7FuU7S1jtD
ssxK6kOxcmyPerlFr3SBb8R1ZUMYf27Jra/Tb3mgx9NfnYekCvt3TG5wd4awvePhhDV1bYuR2xYA
GAa8LSEkswi5Bnqf2rN+CuoDaICpRTqfTuG1Mn6ieZVjo8hMhNkweLh9g9DO+gVp0YBI8h2xo9S+
wOUbekYoSKLxIIs5tmL/aNyAuMuU7oCeUa2y1KY6etDUNmjXQLX8Q+RECeMJ3iRflrnrHDJUo6bL
LMT7vFaoMVmiv8MBevE+oo4vXiIyS4DeXNqR6sQBh3heBnZOJoHGutI+XbUmbQ3oKWtwyTrPmdVj
gXQ2W6+bXyAgQJzhJFBK+Mb6U7qIHp1+Qh+RNQcAuyVCku0aAZNDU3rmqnDMjaPLLlyKXubtVU9B
kW0M0dp+aBWyT2jlr/49JBfsGSWUN5U/n+nx/1KtxJk0NJvk9bMsWXsIy7fMv4VVAzMevdSAsOFk
q8HdiKazpZUVKoVPauM6/NNUw135uDS0QLj0BFGsyIq2ejTHRSaxzZfw9U43QvxcrWD1EG5wzt/n
8K9HlSv4Dyk21O/mlQnSynKXgx7mMno/oCMY5bm5GLgN4vjHybCQV2Mjd/x1vsS6xnu3cEvYKVA3
L6pIq0LJiTv2Ch7z3jhaIGgjV27IvofRu6PnEDE8wdvxnpzlUbAY32vM038Fs59M2cmZkVwSeMGG
81Q1Z7Wcpt86QUc8OpIx2EOqrVvNTIkmXMCxb9OYc4LP7mUfQlZfGIA98GLq1Xat9L4+jR+Gf+H/
K2eTMgHuqswsVcg/bW+w631MWb+1Ukiil2qc7KX6FxP8pwa3GUvdeknfaFWACutKtszdiH0sf+9j
5b0TekJ5eQdR6tUzT2j/3fQIjLEofI+qrRQkp2SSR93sA5ahxOritfZz25X4PwqDTaEA/oYh3Qqm
/eZeryrLw0qgt7x8biFHW4RXtdoy+oaTkvpDScx0ssnIRhJX5dFglhDcqAZ0VpICVTDAUGQmJeZ/
f0vvG1TK+/9fkwJWHrQ1jkOGUGVCweYl4AM/2JA62TpeWE9K1RYt41DayoLHXcR8d92gfpcV5gN1
x0crAVKzQs+OcaB7krFXmh9o2i8V9JZVHvY2WrLEqJpj4S4s9Vdfpf8Vc3HrsALUO0utT/wU5G10
/dD51XJr8vtJqj0403/qJHJkfg49bzhCskp5RI64gkhMtjQwfTVg/dqv0AAzSj2ZqsEerieC1TCj
Gxf5YHq5HeO9KMVc7SOqooWRHARTTamZD1AYd3mInR5ybcpgwzV5LIWQUQFTy82PceHIV0G6ljjw
RUXlK2SLd/aZXVupUR+4+WalJbN3HvPtW9KkqBxDrV1A3vNjXrieEB+55GHYwhQP3IpC80lTMgxn
Lq/Vfo5pT8xg6cx+sAas5vdr75Tn/0rMe1tmSOlR7FRHP4/Of5XsowahFvYICsDeFXiWT6b3cRaY
zkCLrK/nSBUekIaOWjgcllQmawTRXmU7NiGBKJVSRQQyN3w2+J1zFt7aQuou4Sv2UBcf114vB7uy
z6VHe452dZtDVfuCVilEvN5enhueqatmEiuqQ41f1W4l15C2G1/GUpsh8Q/EFv/jZUw0WGTPmdVv
kQ9E2vB+kUIXRUsCsd6chi/Tq0JzGFK0u4KmJ+OJuB/EJQozYxwpo6sId0ImtSUrf7u7J/62dayG
MQDMQT/t6ht18NI3zlkD7z97FqUaGM00K+lb0e5Qq79NhPvZH6n+dCHcBHzkX0oyLCocqNHXVrgv
mtQQHFP9RW9UKgM7szvyxZ43V/fXA4VXr/G4KTKz0T21wRAOsGvPToahFR/sq1OL/svIKlvLouSl
sKAepqOjMiNXY+8igvojsYr4RERTxwsjtNZDrntWXq+Zy+K4FbVeHPpMFgZTkuv3U/ABoM0h47qy
24L7nQrM+4LiKSEopqwa7e+XG0AYH8q3/xSpbYfCvTeKl1QLxYyWgW3IOGUI9n+/pHIxtEr7ToUT
Wj/w7sBhtLJMeoUlx+GLrHkE2CNImxMKh7+AVpwP+Qk4hBXrt31GPdnu7WRGyG0wTH6N67CapKF5
ZRnWKCWgBvwP8YftUZSVSyl/H9eIcieBSRGaYGrLmX+ODScDIax8sdHbqNYmsN0ikX6zioqJPxXY
IQ12rpcpnU4uLW8II3I6Z3KwbT5MgTnERZKH+iBWtbU7RqXsh2VHQcxyhE6KtoSKZPA2H7+UWe7M
klx0WnNSOZV8AryxOqvsSO3MBAcdKCZvAQEZcrRcgD4VEnfsLQQ7eGRHPKpluy8KamYagSNVYhSP
vKeUgAKURf/8W6tghcb/uCgmKOpKdYmczxohBB/TiMm+1Mme/cCiBRZl58Y5Ml1muO94qhk3PKX+
WUiIPbf8ukNLqwGZDvRMiLhFoDsgxgFVJc8yca+VOEy18SLtD5arJT2vPtNRR32TAiBC5nfZzYc3
gI9ijUqDK6KAWMKRGe1bJrsG13zZ6C5wdgBxtJHmzAsfYlafakamwiFy6AAfkfvYYK4MW95ufCwD
dwQKXe8d0RhXEgcOrK76Ljeyfodo++ho993V5mQ6L1p0eEW43AvKdDhLUTkm7apO8wm9kcsRgOh9
BFQU5m5r7EiUpk78hk50nrPycR49X3TuOdad6C99k5iDb/oX8oYdJ/2JSwyZIqXgH5LhRB1GsJsG
hKmFFwlyg9vmFhe54msTyDWvHcmAU7TE1Zbpt4s15dAYbbiNqfrTnRwuKm+u/t77kqCgaKiIvUes
pCjSayltahhujSiSt98HxZ61ozvX1PlvJQh0HZma/lKVj3TABpRyRWAQp5PYQ/Fu8fiAZfo98Xky
Jnj8i27VqB1gUkayrUdZzDCcvtsPAl/RiX4dAQcGpVlk20wwC/vm84ISbtjbDQfWDAAY9V2aXvh3
mmI08MsvScS30q/52ypbra1mHXY5lWtHOWMxj881MBxD4pNr7Hwgzw7jsmXwdNFZLcPlszn0ECi9
xJHn2fKVUvW09TWV0B0pySGc1K91ikrXjH1Yq9oHBT31m80UVqkN0pLm/QRs4bf7MirrUeGZK+Ms
CCfgJdAI1e8SiIefCVGgsFXPGKv3eT12W5mLC1kSi44wsEjmnLm2QHClsm5A2wmrP+qNNmJJCgEE
Q2AUEdeBb9AzH/3m0cwyd2n9xZw+O6Qba8QDIf+2FkfuWKXC6I16DXFdcjScLcuhA0gMcM3Oe/4e
o95ZCL7s7+6Wi5rxzOB/lZnFSYK4efE+S3fPBdGq2kyXLsxsYVzDl6k8Ya8L5aMeSLmkfzgftema
O1YNmI9hwQtwJpNpywo8soc0aqp5pZkrPTy/VWoIljICKN22TDLLcov5X+h72doht6eYzSdTaYyX
oxQQfZvljm0CFDSh/4/+vCB5B7+qab7mPWgjehYGJA8qnZAZeDXymHHaDw6XqCR3/+VCpTbnwWPa
G08XidXbgsgMQzvc1CCa5/77Zgvh2/J6pUQMNmeQY1X0l/xoGG6DFRwK2ll8cuzML5P8QHfcHoRN
7Kw5LqMkHAOlJWyWIOLktx22GWAodMfE4+0HWqJyAk07HeBE7IBYU9G2e2vRlHjDIn7hGaDIkOAE
IwX8t3A7niVtSezFq65+J839XTSnAbmAJ+/uq6wfTC4Oop4/Q0QNjYwyUd2tBfsY/zpOfIHD+MIa
XFkgK0ILJSREcksR0oBzfdCmOHIO6113YAnwV+iJkaZDNgO2ASJK6uG/M/o8ZVBBtTFbxvx7VDQR
4PriMiobbxrPAcw33IudAUJDGHbocUN1FSOyFWXIJAUuP7grjWNP4BEfmm7/6Maq+zPPkrW1iQk1
FkKHnFa7LPhJiZEZhuAvlOP9ueEIVZ9yOmuckTi0r0srFi61fFZocVcdL+ZjZMzy5jDgVGinpaTd
x66/weCIFw0UTLOKiDcxvwnphsR3BqWK69QzqAcYNL3fXUszxhiBvHLITF45b6xfi9qpVuFDQVDS
P8X4ratYT0vxnOud4kPUgAID0gu529mmIUSVIr5bIM3HlsBhQHuKSeJyzBfimbBLOxLYe0FRuBJm
F1WyO65gljOL30+9YwYtP+Bx+D3GtWQ7JRE2zaxxrRppCy1uukRZgmLQ3VmQbxsnLPDcPFlCblOm
fXt7OyNY1aKuH/dL/omxwyjF6xk+F9YrVpFW/w7JEp6AOrpXCtRaNRnTPjmlZ0u2B1pH92LnkzBJ
apnC/T9zALZGeygZyzW8W26GPLDpZWGS0gZNyyd//kquMXMVXOzS6YquzvPga+m15Qj+PXpchBMx
TOiMAoDo1wS7fYunRIgi6ZgCdP+C0qhnMoMfVSbyQhNHpbn3ZTTiQPqlFls9ozH21DlsK5WobRZx
QD4+vIyftc/KturgOSqLNvYisK/r+9+aoKPbqih57WmRYaSXlYCTzZzam1D9XAKXhXzvc+7PqRkm
ndARJYIvWvgi4UZCqZJWxhNwfZe9TntyRKzVRx4GyFCrKSSnP6txXok2IziTWCLBRb/awEzxvqVR
9O2gJX3jxf1vuLagCKbnQqPP+RK4d/dPUU8NsFsOakNROv+vLk/W19jMOv/A5zxOlK00jtR2X/iB
2aW9HUD9HGBctAHgV8mdjICbZy7olfv/MQApaX5SlBoRYHZZe3y/hIfNJ6vdNmv5q+g7OmM8gCRd
HevfPSox7DeW2fdRJlsp3RGkvE47MajR868kdp+Ue4Orya6oZ5FbYG5/wenoincP7BLSSMh+hUGr
CUfiDLMuqFMWyadBRDJYF13bUcbRISY3UvGExEqvsPkVwWsWcw51AINZN8Yv7qrk+dARDRyDv5bE
Lhr4Ys3lYy45h3fx5ueNGRzSfnjdKsa2aiMpXx9BIboMGCW7ZWtRfjwXIg/35HWJ8lqBfe5cg+vM
6Ocf8j5Zk5GxeOFl0U2HgdbrVeut0WqPCR6wfeFMoVr9UffKC7eNTmm/Cn//5YmA9/xXfvsOv8ze
pGoAYufzoxbE1buVKQWVCsYSDfkwYGoDRxbCH3tPFu3KH8212RkiSAx05eAytM9EE6Sy/P7hhIGR
ZiUj0s5T3gLZlBmeE90SMTIaLfkZp1tzS6bj2Vxjtw9JrOKLDAUil5SwdJK6k3xzvbWoOcWokeRy
pgwDGoH/1F6rqsZg16JMmluht6VFUukJfrK88D6qtdljWaDeeewbGuVEUqRCVIlgNbrOhe4rDYn9
tCZp6eAhsC+lw718CcC8oOkLPi7Xy3sGGyn2ggYYp7paqvoOG43hbnK2OtgzRdj+RQLpkLAmdaXF
MskPUhbY/Je+czJIX3cJMAjrnGhfhxL+K7xqR9soejwFgJKCo8BELMKoezNelJ3c51pVmGDe2GyX
d9o8OzvFJBBAevK4IZOdUmYIuSlQzYT5EER3O80EO29lAtysPYMsmZMDXiI1JtTfZ4yBzeIIWcSX
No24TDntSRdQd12gmJ9r/uS31EA4bqvW9kURYME//TbLiY4hzEQd4dwjrFXzzr/9/UnFBfG2l4yg
K88jkSI4teuJQLyihOtg0woT4Dhe+GlGJ5bNGMrqXJTUZJmH6mdlNGdfRI8/t5EGZxQG1NDUtklB
Ojgab8eccCjckCYj+KxCIZIyRYhnV0xUg8Yg54AqkGTG0W/H7cdVU2kd1OMYKoT8FiQZy0qS7Hk9
AfcBZruAXTXebpBrumyCfAetqkuUjucOiq8cj/H9hQXIMvS8XyMNHXPhDp4bYtcvTTPC0+1zc5Gd
FvAGwO2ijhDr+8DS9T0FVJ1ertLV+dQFT3L2CtgEWmPIhonvDsjlKRfhyKZ7CEbiOzVQVjf64Dnp
2hTnvfgshqzR2El46l+OwCbiPWeWo1jyPGVcG/xMrWY8lWyIhP/DB205t0S4h5HutZromogRzIO4
yNB2zmwwF6cEXN+tZ83vfJQCzaLwPYQ4uo4GeZ7DGhlmmHLXHrq9VbVx8NIZoqo7qZc2a7OWFP7d
A/aGhd0ClabVxpT/2RYsPNRYngC/7K69SwDm1rjP0GyTJk5cT6S/hAl9MDm7Xyy5zUVrTkdoNLGL
JTN3x3i+bEUPI8TDvMRzI0ywb14YezatiGqtPTL0x/qN8SzDqtAPm9xeN6FWcdAaRuG6c6r4FKze
PYmst79ji0U94ZE4r+Xinrx6Q38uymHh+DPJxfZWlPywswjL4TvSxoGK6rBfAj4tNBFVe2xhZwJh
eL78YmIOUEWP6k7fzm6JI5nmMusxqtMduJ4VQiS5mcXJBO9cFbZ00zrLepaQj+HkHdExinOXVhqd
WzieoVh1PH85MLT05j+qZt640eEk4JkKfuYwEmOIBpVotHYCu+0MYJx0i1r2UuqyM7fvEyG3aisJ
rXx7aZm6bR9CPVO9P4MvrmE08s5VsLlMdN+Vbu9gIJbVXiWBifITKrOsU9TA0RyjgYziUBAvA4cr
y8U05Iwhwgab4jxNUw9SbSFZD+n/QGKI8wn9HiqyFlcX8jLXeT9TAd9KhSzjmOk3gdnYJ8JZjWky
TIuQoDE6uYQWzu2JglFKqI2H8gbgWCyo4z/EiGypigzPPeTy2dLtAHBtaPe1wh/eDwH1AuAVb/Yq
AyhfHM6PVsuMK9Y3bRbWsMkZCVcCnP8AgciY9IyKIbe0MgdDPlwN84Pr2QD19aW12I14HoVfppPD
wqAu++r8ve+ZU27kbcJtQKFn3Ro7y7D9VUn7BqhDbEfVposz1FEklkf6zJTQAbt1eIMRDtGC471q
oE2fPHljvzOxqs2qwUH3G2Y+0uu0u60LtWMlOFnIh8Ee2ZyziSGvlV788BCDzlUzQCF6qxXHUnR8
I8dWzdgzQjgTFFOfiDzp6aFbCpgdYW0lM9RuCck5DIFcJ3BZ2Yk+CHcWnP5RaX1625gGstQQil31
SGYZ7sm7G8Aj7x++As29Ys+QIfAXF0gQf2e/D7lkxm/w/IYy9GMQ7HTMMIVYcE+lqC500wwjxfq+
VT+eYCjGsNIYOhQ6lI6Cii5Rk25sHeVn6YvbbagEB+Z7LgS/4VuOOIGCDId3pxmHWH8kObtZKiad
enUEGTOF4490YHPUvWJ23KlSZnxc/rngTYrs+IUrgq1CY2GnMboGNG1F7Cw0N/Eu9P9zU44/AmWF
6wh/2QfJ7q0vm1oa5Le/MDoAFwgA13JD4hvs5CzP8jXlPjjdoOymaCMseYe8ruv7gdwPbO8Ug7IF
zg/xwJdG1N/cEDz6BZs/qIWYXTbE6gjl8LvxiQJ1ThIEunvw3kb97scOMjIxBhaRonuYIAxjsNjv
63FvxPW0A3WRk7MFd2huyWj/KOYHQLHZnwYTSl+SoUX6CUkumUDj1JWRTIIczp6RFeyglnrzcS/d
uFj9Vmp9SNjqZuquMGam7wZXvhYXPe/SpMBHFj3Jb7WKV/zOy8yZ3OHsBgkOhcoBdQ3IPDGKyr8e
35TSserWQbDr5N4ASL/k4dq5+16uzJ5h3PjCA04KjNqQqvYvCeUt4rDt2bNsVjOepPNKjoegOXyj
/epf6XbXgysJb9WD/ex6z/gm1yCw33p6CJyVJ/YOQEF/AISvGvIgZoVeQQVHAwWio8bf2LiW2Y2V
Qik8GdM4Ix5+2D4NvW9UbXhJp1uFo2GRBNf65cnum1iwO85HldX7f+M5cXi6FGJy8X3A80y2SPvu
0o/DQD+bqlCVKs+D2qrxMzL3URcsYwtAyMW2GLCAfTV9c+3rUfXyqdQF9kU4Oe1GME3Ce5LOw8di
4OK9pFinrKmis83h2OofeoztdyJMZPFh9W/1TKw/nwTidSs3XYtEjvj1EkzDaZAG8Zlvh7WfanAL
Pb6dpZ560EfZPtcLQSvYHO7P/0ZnEb/bXtuj9jYlL2L6FXHlO/ModZ0w1HMcC6USAD2SDBnrFDFP
oA5sxyLzhG4ASznDm6z07a8Vm8by0E59Uffy2EKNclhCuvgwbYsv4wsRb58A2Mj4UVIleDmyHk2g
UvqRGrj+Pv5Yr1TrUGFYQiZKFkexqBMGvYQvzGjcNT4b3gqFS1JyeMODpHlf2v2CZpDPnq8CX7OC
SdTlXnLPekk8tnvdPk4H+4/dUNi+MkdveDQuivQuGYH4W+hpCNphXT+WFw5gNwOIhI7wZpbKWbd+
EiU2pO2pzBMikIwAcY7j+5e6fuV0+Eu1lajWaUtPLetDro9q5CIzXzUrzmjPOXXCPEVVIu+4SCn3
2u+EV2loSLGRanJpjEVFZUQeaa+P7brjuqkzKFvk2pkgjesKQNsJp4YHp0ERHg+Bk/GsvJ2TCfKs
ihV2XpSkb6i/5mmUrwXnu/qxXWBg7EBSYdDsWrGxwSiPAhfk2gWc8J+gbr2lIB9crMceE2pUQ4l0
9tdxlyvhvUptpcuav/+W/nRcAlKlulCfaT/9sJmccbrHJCAv6LW8okXbqjWWOW+ZOp7C6ZNB/27j
uGES+C9Y/X8ChK0uYpY0nlDES+2l3pqlbYoT3u2cK4Q9bTK+OQQB/h6A5U3Zpe+5Kn7azA8OnAfr
BXjpfJaR4fuoiJcw1qcq+bxUQSFHq2tcTYbwx8SPF1RydncttRkhmOdyQ41M5E1doC5OWWux99AD
C76M4WBF1neNPey/7sMp+UBzAf/tmA8i1eTGb86HTIIpxDTKAtWbSV8HtuGu3oSE+GeXjxwPaBMa
hLeSPTGlFm2ixfj4hzWJ3AmaEbUgdkqKYfSaymUIOVjvNWF5chZt4tov1dGZaK3+r6sEWt19Awbr
TUgLK5l/efyzPQZAbkkv06EF8OJRYNX03aBFWglqRgEgsQBNmhcT4u5PPSa5zw5TKVpg+iZvxdBP
EeKmmUzWsLxj7YYVOyS4yxIWYqXSk0Wov2FLYkwYGZuL2vk5EGfHQ7mly+QOPbyVGnmVRF9KSKgM
8prV4lFtH4fjde5hkjYOBYRAM+yRuLwcEtewU5q2tTXExYX8oZMk0UOsW2UWFyM4D1CwOhgctc80
zI1Aap6Vs39A7Px2DMrOvZuetT+JMLwqCjLpEXe+Hqyeb+TzD7yun8YAxGjxcGA3YREOxhHC6ifn
tfoSRfHRKqpN99VYfN2obVVuTQegQ2isxg+dt50b/nNEmoednFqtK9QPpIMeae3NuuuoP/I/Vy+f
YuF0vuAJRvEUVVjPb56p35kbVq+uCZpRLiT28cTMyZyO5mQd9psgLB+e6SBQmsPG/gqShEgIRemh
GP2dQJK9p02FCU7YxywgZlH+R2wD2DPzucWHDevRMcAKF8TIWOv3SXPETSjq8JPazl/1CaSb4fKp
78faPOBf8EsSMl4x1H5EqCHWl1WyWPWMFay1z2FAdAtgXLwVhR4JuPIfn4mLujvDVLgjj2JAHQk9
QbTQJfvbW/6rDGgU2CfJZwzk2vS2k5eIcv47vwT4utgcLBF0HorFFcVv6T3txJzqKtOObLyOR2uz
st954zCgAryiwp1ehcTVB7+wovdTnSCWOwXUwGzkcTOpe3kPGQSN/7D6uwLFekq51Ry5gEWcfHKq
xgYhzDzlvNJnqfRNARMENHOOkwOkOdEIHNmI7PgVR8ZM5JoX2E8gQilgLJ9/eP6sjHm6rkw3pmV0
bqdf2Mh6x6/MERua/240qu1xWL/TLngnZZ/r2brYRFhLCSv+C33L3yEW9alDgMWd846jDeC8cjOH
0vq8TWo+aM6dSSBw2IjBe0zxlptihZuOSdIiBriTU0G27l2V8Jks+j/SWfxM2jRZK4wRXj4UmLyn
bzGmnPZN8pH4UEDj4+hXZ0t6aMHPuQtbQKryHrBKeYCqMIBu+d3hvMJ7ZqT4c30qb1Y/rsP9NceT
Eacz+bjEA+lN42JvEYCoYkx0bxH9iEOyM2ySBaiYXx6q4ql61ixhZfFDOGJmf8Ej4VES2YJkXyMJ
VbrTeHB/DVTpM9NrI+laEfrm081LJfY0nYiMQvi2n8ClkePTd7vTw0/yYyuWMuHUHCKW9elFq87W
EAYi/V+1td7ySTYgIhrCpwt02aF99PDOo/K4MPxvrbpWCTjhlk2cKWiQo10hA4pvAMYJwxF1+Qb9
OZvjMB2h3LVtBichWJUOLOJM4iplFFzxEfQQ6nNsmSFNEk/wvuynuQCor7elzLPOLkz4hacrQSye
fKMglojZcDamAj+ba0Sa5KSU53fYddWW77bIKabgWUr3bsxvXEfquayyQvDAc73DRNCodMz8+IC/
qkOmroPCTxQehGnZz0EHdzsHdVnALMthTZQnGfWwrTYPUmtBSOycJTlOe4hL4q/3bi/wCoex/Tuc
/Z9rQuNi03l8uSPhVe/EqLn7L1TEMgMxKLtF0G4rfxJ4wQzlwbhinxv5AjMonjBDcvUOine76x9i
kx4HUEn2phB3DrU6Iml7OMTc18AffqmOr5mL/FF2XnSLWI39pjMy++fvXGvX9Q+hZNhShRnKAKBT
Ugp7mhpM9IJvON3bq265KnBeqpE85zJSd7qPmNRRxbcO6g7VZPRVqkI/pyToLnp1fouQ3oDb1YHb
5KNX/ARvx8Pb05j4ed4V5O73XrTpKMfDVHK3cPlZMS5bMS8nSMtUxI3iFspsl+tGKgoZhbjJOeT5
m4XQQv0lGCDLd/tehIaFuHIfMapnua0I20t0838IMk8LDJsWoWeQT8pUFmvCdjgyI21v4HktaWNb
7iH3WkFf8XvJUFxygoA+p7M7ko1RiNfTc/piWvf7Cvczvn0VJpA8LMPJhN2b1S2UCKI3QCLnVpem
YqWEAsFOUxURPeg6F1397GMo5Vs5YMziOJ/LJ2UgRHv69IoAi4L5qBolPg5uXwqbmufhi9BTNGha
qgP2uE5Z+UdFapn6NbGXe6iNG0Bm95iahRjEB61yDtGXG3zggSG+thHgul2hrEVBZC4bybGH8G6J
7YjENQQRJYsucV/D4d8JQY7MlOIe+TyRSbo24mGwtDV5rxngpC+9uM6yy+ZkyIv4onPRbNE5PvUS
tCTNZFilpH+CFcvoJrITv6JbOhehy96mz5OwhGVaOV5N7NNq1csdVs614ZbwALx9lkGhnrZFJR02
mw1L3t5hhMFQL1CpbT8MRbWwhXyGcxjLQOeBQmydmfnmL18BDOkfgtlzW4YZMCAskJj9SzdQuJiR
20/DHV+g1cKcaUqUT7HJcL/ZDxoe5KwDenLR5z9b0gPeN5WXcQNXlDzZMqz7tKYTQxDVWDo2/C0G
lMmwnsCqN/cmAxvouQfsoi8X3mEF4rEVDvW4IzV8wB1wANvBm0B9Kf6wWkarhWnZS3L8BF3Gbd43
FgtRbzaHnhC3IwW0WH058IaRjNThXTwxZAQLtSL7LNkBlqOM2K2FgsGBKqlGaEhiNE2g4a0V1WMN
c6yQHxmQ4cp6s+au7uiOOZh5AgbfMr1EXqMWfyFLw6Dk/8wcU41xN0os5nlFg/Ope8TzUjXzxTSu
gv7Z+oqazA4PwnESPbv1KJCMS/wzQUz0XQaFASMHCAH45bqlzNdVwrLtL+ZrGnCXUxMl4Om7ZUxk
ONEnP8ZRVl4Q6+ioknw2MHYoVpTZvKgdhYrE3wgEsg2TT8oZ6QP5YeRIaXhBc8I3kRisky1L3/q1
Eclpr5oVbM1nVX9VLnWotOOkoUu8p4fPXfdRwvr5I667mMchu18N1pj7i0dkAN+qJi7S63q/nBZQ
RHDdbZqSy7D9ImOI1LjAB7zQYBmCqHrk6VW48SBiZr7O0MEDEthKJCViD0thWAlHGEjRzXObaQyi
wKXD9dAodb0hR+aL+VbaWA1TIT5Jx4/+TeZjK2FuE3MeLpIk6ZopeEl8/nomas5llK8Bi9WbvJSc
BlnUeqG+gqMlZFwUMoI7IoD97cCfVtXNYxZKdSHDcemetdfPJhk6EbVVKSSsaqtE8v/kXokLwapH
ZgHChjDCgWdWx0/tQKIKXGoh/yzFqNuDLz3z2fFp8hn7TjcHlDp7j4DhDOCVK63cRRf69ooGnFFP
6NmCDY4IFXoZU879Q0sTGD087l/vjLjdq5p45r3C5oDdklcvcyhuDUUAP+u3xPa8FyUebc8HdeQt
BnABG6f2X0WbZ9dsG6SKL/eO+TyGvXkQtCT/HmCbNNd/GWUzz8VU09cweXriu+QJDpD/dU7pT35m
Hctaasbf+bco2W01T9rWAku4t6sD0j5ziRaHZ241swVMdwZDTirOyx8eRnsqQkhM6MigdQR1MD8X
J0K8+7lhePfYMU7GSivrin2lzXDsRfV+F5qNPfqMA2jZdMclVklmfY8Pqpusw09v7iMk6UdphgDd
8+7yoO7ctTnOeYL5vWQGxYPsqGkPUlniw5qXa73r6iYuad+vu0GvVNLkIUyHLzlSVQdzV3RQwePP
MZtPWeoi108J1gdtUAAArqFd/ESybtr/sZ50ljp9EgjIKE6IUFgxvCO6jD5xyK7C7w6wBr+Q988d
te9VShrnXJeKk7aHQoJeG/5BvC/4o3PVIsccgzLdwtweAP77RNsrfVwUqLtjQNVWQiTEeyAX3xk8
OBgjlCOhCaH2UZ5zA7KmP/LqMYp9YJEvbaySLdeuBJAX9LrkOnZ0G+AlQJSGCXpPUtYnkffsmreN
XLuVA7VmmVIoqmeKgpeqR0sTIwEehD94dqdJRi95y3yVumNs1vnHH1UEs+ueD9fMOuk0xlwJql8p
0dicQvoK4MeSJTGaZ1F+5/KGAsUGbZBPhpYE2FYR9IPVNT5EIU5nPxgA46M8J0WBzFs9ZYW9otGB
uCLAVXzQkoWsYQ+1/9RJ6IPUAlK1RdO2op74HBQT3TDOtpHRAdj+j/btrZ+iTj6FxhJVZMZhLCE9
9Knub+k3vOJCMKM9V2qYOYJMLB0fYX3UAv8UlCjo7GOX/0AoknXfXndHWng61eDm7Q8M7wsWlJTC
dxyeqUs6/2h3Lv57exgXIEzULqw+vxX81d+KfdclhhiLLpfpXvMgNyttxajNyjHzN3ZlRS8fMjOu
BKKnS58V7sDI1f0EB9F6MkzLwEu0Iyu2xcCvQKNLnl9aJTv1/g0+kQwM8fkYcWgQsCIeEAnLALm3
fRlCQRWQOmUVyowHLobnsuK7zB54nHAb+Yj6Bm6g2Djw0WAVlMYT3R4XxSGuBP5ZS4LSTDnExyWH
LUoJsWizIeAEyrIbxnZjgvJbXI2cyNzfBsZa4+/YmrdFtz6vJQaPnQeuw5myHd+rIViVywb7Q3g0
8E0BcBMH58N1ZcvMaa3LPahm3OcuwAaah2uOCFogK/QLt4NgEybCgPz7rKFjUYk0EOEwQODzzX9T
alRU9QVOc0jDFUIicGy+ozItgFLk88Oht9SJDezqgXNZG69XbJLRdynNq1bAkgoD0x4jQ72JdmW/
sIto9v77BeBRr9jZZcqiy/Yq06U7I1YQmzhwCUK3AsaToGv5vF3Wt6kuJxKgebBxjgsZJcemd5KL
Y4w/Oeh1JhcgaAfRkt4N78xnOZfBjmYUJsiFpa0d3Drctbt081mr9bgqziAQzrid45oV18iBeCfr
q9Xle8quUm2j74rjDzPctyhsl4jXX4LmdDPtorrjESeedi2TpDggVm94ZD6wpIqj32b4SOsXcAiK
Xt79LP26/EpXgXj8+Vc3lMCoJ5Cegk5QUPZRBDSY11ffHunk69oJh8NM4cA0L+yZ0jK2e9bKVQW1
nb61CC4lGKmPZ6foY5F6nPiKidOlD5WQV6Jhh3ldRG8bLjNu1YBLKmKBjaSVnamUN9G8YxOIoU5I
52AMKPUbixs8z8fvIyr3kQ3w+mJXm5Nn3NlsBGvqDn1yQZ4KiLfN/PRlE28+dgMIk40HgrRz699l
1nSvUKqPau3XYhr6L6H8xwyy2Y81Ka9MmsWWaB1pK17k9YwFkozjCWPnhhaFXq0e71MJA75IvI97
O01iPXXEmHHYjoaxdXfLMB4f8VeMK8zz/RBUGLD/XVhlrKLt9vRd0xmI8HroeDhGGRZmtISwVcfV
Nvw6d0cCT2NPe5y5//q3uwD8ri1KQvTnLticTpS+BlpE3JR68tJ4aywalLI4dYH9wPLdX0BvtoQt
EB6+BBku2Wt1lQBOr9oJWrjWr66SSZj3G0nfrzINrzXtHKoh07CQx08q4LYsW0r1CD3zrlX9fjZp
3oxXg2qxKFXHZytDUuFEwJgFjwsVx4BPujtHRZVGlti/AcS5kBJnydgXKCmrIJi6nfX1vF4M0wVe
tt0nfIZM04lj29ILWKs5uV1/YVkU3ZPlfRKqja8FDEtaHN3HNRR18hYCS6UwoAk6Ck32cjvbP+sS
4+yrLNVHkF+nx7FCD5myqZQKSGUROHUvqro9eH24cd74T7Z/A7Z1yiAKEW8ceYmr16FJzraOurwA
TUEBlddxSdYn4+V5sET5ZIumqu3INhzxSi/ebZpu21a1K95JCeG0+yTfAt/NOWkh8GBUobBKpcf0
7aK/4lb3TvWYW2hquMKwCm/aEp9BZ4DfEwDHA5eoZGAcasauSSvztfSiH3DCtc2B7RBNwTbWpvJk
EDSdFpV6375eitJRhu7oBsG+zx+dKHWYF0edNgksX38I5FhXfh3n2n3WPjWGD8zWl5yBra5MgHOO
cmr/KoaRb+yqO0wTKM4jU5cseX0Um9EQmOlojQrBwOQbuUpzqdHhEIn4IqIp+FK4Syd4fFss7BP4
Q1zBYrGdpQXqRauBT8k2tXdDtWR5dSz7/u2MJ/nmkniM42oeL0o8qoAtf7C3rzgx6hBIm3s1mAMm
UYd+ay3Z7glji5sRYGY9sFC8lr6lLczNzlRmnukRbgIHYpIS5HvSzCoGAl2RVp1yU4yw0hog2wcC
MXV3VQnTu9C7Fd6SgphlYUGOlb7KYR4qIVNyFvFwbmzgNlHX9axpXs52f5otPsuchAVDlrTjSECA
Vkn8ne8rHrGsvC7MucxvCQCRDu4HCKZFev5mkG1GrdIxFJI+5GsrSOF5T/ETeuqqXlnx538rjly6
lB1WzbXlfrU7KjrVW/2qHj/WmNguILoBGV6heW1ulif62iDJ0ySZaxJQJTeHbLWvoTgTVx6/E171
T7lLHmui6/R+1VTyoCiRJH2KySN0NyBOMHEKUYlHwRQwOqUplHbpMsti77DMFQ5IrGduh+bHyct6
PiIGM0UXtPnSnuFFWSIApcHw2RmBEnzW37D2QwkcvizcMy7Yk82WjydtZDn/syobiFalY9Arn7+1
ydht3ZU4eq7uhOjFMJr+j6BXKYdaw4urzuRf5CDElr3Ns4tKC/olHGqedXNQGDfQzbsyYuw4D2ib
eeVx3Em5k6P51prJYSgo4kUhJOBK0aq90gFKYuDI8UJyYENYvY8h1rM5xtQ4qVMiAeKaYPTYU2xE
FUCu9TCt/gD3GA843x6cxOtClEPJfRcc2GXw4HYy1rJg5eFE0bDTRfAfrjLXStvcCzD3Z4a7uGAt
1Qp7Ol4PBETjMAYzxrsQI3eYnjinh+AFz2hebN7VduDSoFFZbC1f/VBFq17LyGCklO/ZF+J6TOYE
p5u7Q4Dxia7s78MyXRGv1fZIwwAYyZ9TFuVKJ1cqKm4PG9RbC24oUyBip4T7Gr2ZQy5OLA78uk7O
hrzBQ/scBgPJMDF5z4gDmPGvG7KPYv3LWZGxCNio30XBTHHvpcafKzsIp/x+u5vIl1DJ/36FIsD1
4BvP5V1bTVBBSjOBfcdrj66hPj2ZQNokAjSYNGqHZi/0azLQrTStZD/utCNN1mrYObt3v77+8aap
6f7Ul9Wt81s+vdLBHr3/x0LSoATB6St9TIqBL2yPCoydl9AUmFSNYx2jIhudEfTofCJ3agObyO2k
oI1AqfhJC3dF42X4iisAn3VHNDPWy9yCQkccDn168uHoaYjoCkPo1Cusr3MbR3wALzJMC78qj4eT
B9cSilxf1XaSgs2is586/NJH7dXwwOwE5rEYBiKZTBoQNEUIARx2C/1ESxTowzV77UvdjXYkD0RS
i21++nxKPAWkQrWe4IVJphUx84nYG+sFo9Ox9jJGMNnjNQoWKHNWZztWd7KFy2fCHutuLLJrl2vv
GFnnTj9Ww4vdIgy4Cw5L47iFMleLMwZloQf9IvWmLbgUoLA0v/YULtjedit/tuq8idDSJ97/ZJcG
70WtbQAdUzuGdP3ReGFr1cioqWc7qHoHj1yalR69Tf/2XEVTRQtsYzL38U6vAPIy0+Y4Dq6OVK3+
M2V1wWvMTWd7afJCRh5f6FVHg+rqRvzz4l8oujdtXsUUL6hIthEocUrwNcQ09L+mAu5u4FzLgDws
9ZqfZpJ2yGXMOaL7Onp2YPkrt0bCKv6TNhgViq48ATLoBkCrxRUQOm5pDmYT5mQhjVtRfW32ZEWW
fLf5GTRXEt+55B7jfTxYlHhdLUB2S4wvzZs880ySn8Ghz5giJqLRvUHdgoN3d++7zFdEYj8tjSV0
0ZjNKnqJwrAjOn04NOtNcRGPOdSVgHUr/EFVK3ooTtCliNRBcop/zU7MmKeMNswmC0nWDpNvPkci
BE8a+NGx4AFlqIIp3SVGgfj2NUM8a8qcn/C/VwtvfzmGUJhoqeG6jr+XuGGVBCg4M1w2OP/Pu/SV
lwP9hKdGa+JKsC+EAoWpuek/UwpqAqdcy7q5KXnw9DOlRbnbb7jkkznJfx/n0W/N6R6y6DT3wpS9
E/rn138+KPzUQEeG8DXY4R4DjvG2WWdKQmMYo67uzPVC2Mt+Of2BiuFnXWhUGZ0bO5Vvr53vF1Kv
5tnLk1DQEK/JneK9kJ+/C5oP5ixzzHCgZuR3mbuy65Y1jHk6OkpVg9dOe3VNgYUeK0YfAZlVlhlc
M6QpQVMsdr1Yn1i7kppz9mUEEdrILwlKgL6Bwy6ju85GZl65l5FuxNTEGjqcZsvgq0uZg5XEGU/l
FT0B6F0JirgNawzFc1CuEa0rrVgRVrLKLCypVgkZNPcLqIdcNxLpveSYUe5V2/KLHOakumS8NDHg
bAy0P4a48UDyhvUrce2S8Epqvo2AU/L061ZdoY3LJRAZ4Oyw6Q07XvrORlwAxTbiGW6fMiI9aqky
wuKSei7r0X0Jn8bt7fGxk9tbD/kTj5DFg9vhUwq81lubRJxv/ekRNI0JNnqZ1se65zVqbNBJQji4
X2+Wui0EEDHzOKaNuWDSRUPpuN8ZI2dHZlzvXhsGtnKAL/95DExw5S4o3mqWpJ/ZM3ue47wBYJCf
DViNHjMuM8yzxNLoq8fvLN4W2OMfRC8RJKot2UQR4xkRewfXeDvdYgZrW2k9rAEqO3poYWyB7GRP
ONyMAx/BdGdHqcl9H7N1EJZBV48ns5OoAWcNk/yC+GiI2ZnKNSeLni2kGjYNhFIv8IYkPyqkWaKQ
7R9YuxFAyVq3rrFW57MVnAOVbCDCPLQKcjqGN2zNVNr5Qc0XExf6b4TgMFA+G2CN96YfCq4zWd5F
CbDnRdDs4Uu5lLmVY9ezcJVez08DebJxhmx8fQhE4RfuFuaXpVpkjdFx01SHh0NWu9BfVreIXn9/
SMq7QyT698B/E6999phJmQ2i8l/AHcM5lvYWoaKFOmxr27xzr1jZEdF/8SPHRPrK50TjcaRR2qHZ
M0pu18bR2qVM90pl9ShDZycSpElvAXB5JjB4co7Sf3ZTyAcpf0Ym9yfP3rqJDsMfP34xcI6dm+CL
E50Gz28IRxVxPn1ndiRzFm6S+vQf2ypo4KftExDXBc31GY7d6OYEwIhnPRpKKN2Sim5tyZwE38gY
F8XPEzBw+I7Vti29UyoCIagouzq767cDOXSCG8r5/U7oUrEEAPSpv/OwNOoUesUo4nEhIUL/Lvv0
c9fxL2zmcQJg3brKOjqKKnr3e6hY21TrE/jZC8rtpXZoVOXTgZXOdc0sFso0+jrYpvPYp51I46UR
fXDSPt7X1auWBEDe+KCH3+7kub+0oACIX8Ni2jY87LXNDRsoudUOa3KaDq4LGQL1Ea5C3vPDycLR
OabKmMGvCXPyWz1WqGIdioVLWqRWwux1kLmmKU1fUK9/Qwm7ylqMcnCrRFO9bMNRicSooI23rikz
Vald4Nf+P5Da01c1XLRdEuqnTrfEASLzv5I5sB7WZW/09YdU0lofIxlPmdepY4w1k1zJlenG2KqT
XFRkuhmrsNcCSWZeD+4TRtO8rSKWQGukP+1Z46coZ7G/Hmb1Rzrvb4qmHylBfaop49mq0RmKiWg4
geiCzdErEta38XAsZTUCTJIjTTjjSjWI4wdbiA3Fr2x44y8ccAnKDhMHwsrSJXmAV8Dq6Z9lnS2J
rx0OeYSBWX11LtrsLB8EPTJO3V8LNw87wuTXsHf/NF33o5WyIdJsUKJG7G1QpdeneT/vHbaQzO2W
r2FeE52j2ID4MrL0hzaQL18WkX7NR2934mr5pKym5QjEYY4FFvM7bpohENr6EugqlmV5y83lPcLL
N/iplwAgNtchIMyZFW1lkNTfZa7gi7kBovkxIrLoK/G25Gowevr+ID/jW87y0RbEr9itueHpCiTE
0MkP9bIem3mVJJDF9fqa3wscLMGthOos7Mb8CXMiYq3u8E/ckCSXZAEXyJcjy8Kg4zNcTPrR4Rmo
0BTH28bDDE+nmin2OUqwME4O5d4v1oq5jugu6dtPBWM1dLJD/qXTsmbZGIF3nGwRzvxA81RUQ4EP
uF2UDdLKIOVtoABCLccZ1yIuBK55S6ytOwJeogIUjc+Y3ZdRSM265XCk7TkouHAvHCOVaRfGY1tY
LYsavK/0dWTTmW/a3QQG8x2e73PeIseNNoyAalpe1HfY+09uybfy8tdwp4rsh29kIlCDyxc1QPIF
1AIsGoSLADchU/jYpmcs1UZVuyIQhy7bv5BdSdX1l4C9I2ZD0gUOxWXFnKIpENX42EAxfWcZPM75
Xk9DQ1a+SaKQfo+wnMsP4YkOiSXrThfpJcMshVdCYadFXAsvWEAkk9863MQZbt4+OqjsXIVv6RxM
XTr6IdyxYFq9iWgNynElTrFq56Gt7k4Z2Ki2+a4B8qIphn4MMC7PdXhwbG6+XtEOWiprQifOAzow
UMRJPXwMlENzr/+DWrv6UxwrkiDsKkqS5Hpv/zqURt7o/Bttc6EnD7e+nw8Ry39UdODOcHdScyef
LI0LJ7iHmFuLUygQrrflsmyIxqKtiJapVrOgVYyp1gVKYIwtK39jjeB+UDFuNP9CySJ5TiyT5mtd
G9JMOp/cdHKJaeHhXBKSx195a84ZM2taXyBMveDoHypNt+JEFkJyWO6SaLLwTJf4kK0yUIgvcNKs
q29Dc+OsBJpXmOhvRgduYkQlPRmxhu+Bak4gFlCGJxvzUZX1VmawGGfOaysJEA/wOAGY9Mo/G6dU
lcWdJuEVZjlgOcmgeTf+5Pha59XLVwjMKEQr44ERCEHw5UpyTOSXSDwSlYjAGeg0r3fpx8ESSE+U
FbMHAqNokMzdYyKN9BRzqvymJLg9ZrZ7Jfqvccsrtd5Mtd2t54lwuJ/IC/BBLfF4mUDU4vcd9oJn
E/QJge5WuF38tB/UtqluqY7H68PIOVMi39Fg0cKlMljfztOk2D484fbx43+JZb8LdHepvauL/8FK
x4Fsv70QCLXB47pjMvqJWsvpAT9qSsPF2nYHRjrX4Pxd2M51aUhEgwY8rp7gGMF0/rzgVMHiFQri
rhNvhCjpsmHRnTi1fcV0TIYZCc1xR40zStQmkFwyohgfyMiSsNKwzoI4XrU0kAy2G9rr784pDXbt
7B/UTtg4KZwwm8rAZ5x+26LdxVDsMig11CPFgDwCkepoJIEVwY20D9hCsd+0LXM5fZLn7QwBKAiG
8xqyNtzUQzmu1LyJCJUPDO6vemtj+7+kM8DTSHObMSRwvaHm2UF3fV+PY+qUc1tXOMGJyPcCTl37
1C+Xby0imJFWmNzB9tSmKYgiDCtcFd4yX0Tgaa1WRavk57cV+CnpxCmR1+VV4kPMWFDs3gc5ZPhc
Ms/69hIquBlYRhCv5AfGCDHnG5JXhH90j6kOpsz8kyQ9VuIq79pelWadLV54MoPRUr55diQZ9nOs
fXeuHJLEebPeqdjFy80zaA1z/3BAgIxq3MyN3Wpg92HJ6CSg5fs79WPYUip9+HX8GuDWiNDylDrT
cfezP2wYp0o+h9iHmFpeOvvttV8umeY9xa8a3u5PDkGnUDskNsTACIeORbYpy5/aRZ1idmtCvnYO
8SEQNAbOoY5tUHAISoe5Uz1rDwbORt5STQBuJn23/+rQ15Ot5BlnIAHpdKgEZAaNLmpXjNAV/LzS
NFiTFsT8bEn0gM3QhXCaLkFfK9GKtXCZqy35ROeM4F0d9JHIZqugU1a2fQvTPYfzhUwnm5mrpMgn
V3e9xKG4zbIMvd6dPdfr7VD2h80jClzPQJN2mVVRdV2GBKA4/g2iFryziLLUABKIXM3tHLpge4v7
YX99hy+0R5T+3MS/rt64bcb5o4HJaDwQ1WcLCRDgnauzd4Itikn5i2XTi44kQ9dix1OHblUTYJIz
sJAnX+6r9WFN7CJXMp7Dc5cWvIo+nGWnvGxkZvvEzx22Qq6oyFMD/OHd0x3RvdMNDJESTCA6hTQX
VRwSosTaS9xoqZ4g7vP6E7NSe708uIhPI660ZJLY+TCTZnai1JkedozgqIIZ9Rgp0MeJhRrAiYlT
gXJY7Eekwb7g1gDIWcfCR66mAHHjXeuF2LC8RUmf0JerLG1t9dE/mQLYp0/4UF5t4p2pCY2sFu1u
JrW368x/iaYfutV3juI0KyUHlJe3H+XqBV+sEgNbKLN+VGS3amiRuoNBIv6cslLclFdLT+bhZ8Uv
yxLURefpNNGUzCxZR0laYJGJFiyzspGHEpI1sLaYZFvIRhFtoK1+X7ob2nCeBSdL/AnxEjCJBuOQ
lY9nRpd0LWisbB/DKnPHooNYp8wjxMouMN8m+/EUndtShUZDsuMqJHLG1VVJzdaJ1Vqem1AA8t+x
Sj9SFQ0rBDk2lEhqjOXCzi09uAmMSsOII3F46njSRgy0aLrVNHtKB1XE8n3URXgD1ixaSiPURx7W
F5+T3aBWtjvS4AS4nL5P59CUWWcqkwBKSneCCVPm5dUcgBGI3ac9YsRGL6r+Ei214MFdHPwE8hX8
/IiystaDeCfwgcI0UGYFwE7xufhtgdxq+CuMpS4x+fTi+TJZoBV6S7BSnUgVoHapcp9x2o3mFjgq
loyNaEboYDXOPGkHqYQMpvbJleGht3FEjFXbB5juJAyR5z9UU//9qJZOfo38ulnKw5ON9gwYbWmC
nxznKp5T3QawzMPqiQPcXz+AvCtrOQajTDa77inZgc3h+cFRpVSrJNLrJC5MjA+Xh7ZQwVI7CU/G
sOELeHVciAO8IPVhFGY61XVyt9eOySbgFtEJPoxngM/ei/OUeITP9oCAMe9n8xKD6AvSABqmIS20
E4HuEun+9Bl0sJezuwjBC0ALk9+nUB0+J/OEF5k3EoSYlw6LiW12TuhArGmUoeAGZuvwOPy5Pw9Q
CayEPVE7fAdfmMVBys4poGzFYxuhZuq28thY2/ZuqtIHwcuArGLeFuIyFTZSGpk/cJTaNLt0OIoz
olnFdFZ21aImBD0R/CjPXQAkUyWXT6DoVgKRJ6amYqf5AxubhBXpErZ7PBYjKII1vD41T6cLU/ic
VdwVIyqRQ2iJ/d8jdI2wOqJd0O9XBSj3N9ou7SmgOspfLSLvQGaIDZ+fDd0whOaikyGi5rstl65f
gS80NgV0WSH7NFnoNC9hu9k/180BwRhYtoXoHIQtDD2F78m+muE2YOZ17RPWZ7cVriyGhWBJDH3A
Cgks65gUcGsvJDd0AtC3p7vJQIwN4QRta4qcoVGuBt1pWqxEuDbTFRCVW8rMssThkq6HnwbbPV9z
clFHtS0jU2ykwtHIXIF50pjGXmyFvuMb4Ec8l4+skV5tvA4m3cLxA6BX8ehRpv9lS4wKhwHyfqvN
+OxBZu2j300TLc6fx1ymwTvR3FFpNBWgH9weYYdhsNWVQvUumFN0GARZOtzCeI1tjLuT87ie2kXj
5CM52o3EIhmdORsAtbA0t/WQQONmklOMYDh6iEzCZwCo+s1AxoDf7MjtYQFRgb6vOQ0SMuvFh845
EFJlO1pHPNsdwq7PvFSxgs+qqJQuJAV4vKIiiZvIIOo9StetMSdSIVZVVrPKG6lXJMqsoLpMKxWP
I0LsYYljS6llEC/ScnuNNci0JIUbnjQk6+utALbG1ez1BfHxXFL/ggQJjtXTTthB+yxsPb1QwR00
pnGGVbNnG5m1bK7P7h9mRsC1FYA/4Inrupp+H3b1ODC+lvFzzUGMHl5MbHi+B7ik8XEirNGejkT0
6DMVysECbByRD2zdFzggR64ii/C5JKTqnaGXelnpZqhor+QrJMNJ4TNWUpDHaM1wcqEI/hqQ/6tI
5oSrDfwAJ10nZ6SKm3crWm/38NWAmoql6LypAn5+i77T7JmgDTxK4uC3mFYP/PRqLk8qqGO7AQdR
VWYyP7kkOPPVOiCSLcoS84vmKTkWB0dhi1Lw9r+XF0C3oCixutggiik7GMkigH8UyAZd5PTK5R3q
hupYUPmr6cDyU5gBvY1Q6GXMQL7gat7RvX4JRz3SwGwUfOgKIyWebCL/sbmHQbw0RR5jh0Qon2lx
SJneijQi7GlJWMq1k2E6Jv2/vmlz1YQWrg597leKKcT+P6nMEzJLVfYbj5nblcnr/4Sa4sx5abqP
V3L8/vvKpH7rdjtlbapCNtfZKTzxHKonjP1qTNJiz/n8flxpET4JbRu1FKapT9Tl4kzDwNZj9LvW
AClxrO9WG8u3wLycuC/7TBhr+r1Wu/cXRi3CgaeR2BZEgcWcIgH+uQWf9hJLD6Rmx5LJdNnKGu7j
RbUtZ2EXdu1EGD4ZCqZ7sHiuBi5I85AFqq+Q9/dQE7eXNRWgn2wTE7KbO/Qr48ckF8/PGWGVLoH4
LjeKqaBk4d1fRw3XxoJsJvTIF8s761+VIEnxJpLibcPICsRfgvceVa6106XWZsRD6Def2RZZUPke
mrtKg9/mxER4jz05lCY5sr3yNzblVGaPP5kmHwgu+6kBRZ2u37AqEGyjOfDy65n60Umun2/89SCR
smNlviAMWUPrmi2JPu6FZe/VaVNMEDhYi4mZ0LWOfaggz9gIkugQuFhkZKJjUHR/sVq9k16mWdk+
M4JqcoU1aZtY7uRPlpz3uw9oS6LrwjhESFteQpQ/fAefgvkMxsBGudnsBU2UB7M+3uBqRzLPNE14
1ayctBUswaBznYq3WRGkqojqAd1GLCaW/6S7VHj0d5a4o+sdQFpnMvL5YlqJoxU++1o8ewlgUqVF
+qIsxMPmENsFRmHnCoTwy/HoO5DQcaLWs4I5FxioqE41AzCftGk/5/1tAj2B1IZAXS+yvG4UmlnR
AkyyKllnAZVtIS+eAUmPoIzcklvvEj3spdqIetyQkd5wowfaIzynyzzj9wentoMaz7Hg3YsLdO4T
VLr5IRdMRZodLgOGlyEN5mwk1ONnkuCtkBjFqdAAO6J6oxvY5j4ebZvb7WCiv/FDEsYykOJQ2SuL
lAvt0SeMglpFwfOiIlDWVM+xEAOz5BrMhqq+U3vmudrWUNDyryk876+stUCLeJ1bhazoiuhb6X7u
qxogscIdJRMOqxVxVoDVO2Z7xTNrn320OL8+OAGPyLLPcicMzNQMyVignGnhI0ybnkMvjui188Co
b03yuZGAN7njJUPgJipWeDOyJOT6gYT9FRFVGw5EQjLm/xNoMgYR8CZmADIrxwLTuNuUUI+1mkrT
tpBNNuNOm0TSLO132UyPzIVL28uUUmAkLFoLdQjO2w18PHxRWZYPB2oqKQnt7q/5Tq9ipLFAVvpy
LPpqPePthxPPI5v6W2tVQDh3ZcACDEb7HAorZW/5FkGSBHqfLqBFX6iFLfFv1Ztk03Z8JkoLLXGk
MsBHAzFXDxIcXfF8QGV2nHH+TcoJy/MIRzOfyC1737Sm/zYOF8ASZ/ha3lCsEIA+qbe1NfbSgXS6
wMsGti7sRZ3G5kJsv5rdvg6tVTfXBIp6T0XBrtpIjbySo67RjCad0friAe9FqrKvppaVbHyqRdLP
yHXuDxDzpMH04D0QD0j5VozOUalX35YPB8lnVyYG8u7+/rLQM3KE4mOYFk2ZzD9/WTIRCOK9nH0K
zq5anm8EkFbJIlGSJYZ3BNrMsILyMbY8Tmmwhen41YdFlm0TPETQj0Fq/fn9sfCIJa4Wo4TDgvG0
cB8q/HZQj9E38f9UlzvrYlPWY2tMla+OqIDxwC6RHI48nyzDgunm4H3JJPYPNLKJBwrN3mIhLDhh
wCQDZrcVFrOM0iTAx10Mr3rll1hZwvPhClInM+mzzhSofypgQqr7FoGH3I5MNJlNO62d3QDPMjT1
UCwq8fu3jMxH7YOqah0nZOQKQby70UzmjH8pcorn/w1b+D4Hkp7TxbtLSfYOLokkG2Arsd6z4Iac
smViDQxkCJmOTxl+TP/XYWtEeQRWdNffQELdSAKi7KlgRpprsMvWTY7PGAHRv9+ZwqSC+zfcy900
VtSoRr8nkfEp6hMNRRxHa1+vmwWd4mw+uRzzXwJb/dsiCgO8wU5x4gnEwoEBF3VUz9/JLwFQ8cwk
jan2OOgpb6Dh2sHafjAuqfIuIjkDTJ3ZZu2U76VIvZf/UW+hf+DBva4s/9SoxVhRrfZLeGQTO36h
tvvMhGzaSlh2YdjT42G/YAVXjt5WdiB2HKVqrq4BhaAE0tvL0pExwIVHJi2pNLHxMWq6B37bKIvw
Ewd3l6eVtStOMS9dgKTW4wlimP6Fl7qT9wmCawct7QhXwZ+MxigNkVA28NTOjc3N0kupqUApu4SE
oCY23B0CxN97n/b4pDg2iXqwp1ssxjPNuusjCMwg0DGgDWQzTrlCQ3eQLE16GD66F5HwndkA4Udy
ns2gbMPapDMchcB7knpMRY4oBntTL3bIJzNf5nwxeZ0hE+rZOpGUajZzq3FpfrKqo2RnfeFEjbxU
cQRw3DGMVPVZg67B7RM3e9BDtRgWYjubFAUl/pDY21Vh6VD+gRTxnF3TkWDO3m7HzAOruJkxUR3y
MbLYreszmuIAgcnsmy3oyYm2eIIf2gDvWFmyAFfTnDjb6y1HkBRNYIqoKZhc+eL1XttQmvtPuyb6
EKi12SYhyMl5t4WrT6WxU9byQrXkiuhnrrHgK9/nyVEKujnZ3FZCKUD7D62eGcmKKhWlqD27RRYm
InWAdYsNW0kSKwhtFdpjbCq3EFOFR5tOFDUcmPbuU45HfkaHtK1A+SCuxmBTVuWWmHKVxEJWqEQL
JPItLFCABfD+HJUwjc4hV4b5T0dT4iq5KeunOdH0wd/y9n3aG/BE7fiz7pOMx2BkPYCP3n2d6qSR
T8uKUyZyr2wdYZdk39wDMQ6BnxheZpjMOS9dzMKZtFSSkhu4KAqtUN8YqGFYkIo+h0TmbvO+MzqU
crR7EagZ61TtE6vELUQF47e6bfRuLJ3qItgq1HvzfhhMjMt8BRbmcuL1MwtSSLbjbhD7aSr3ya9I
bEa0vVsbZ5Zx7bFX41UvreNbWeJe8EiOmg0FyGw6vxw/M0086UE8hYHEq8xKun3KRdCK9SqoMf//
vdrJ4XAz7aOlAd3KMHnkmw4YAmNb8pdoQGYMnwqPMtcXOCFfnKNwD//xtR0UHFiqO4fInCRfGTD/
QiTu2H/kYdp88j5UyYOz3Bc1Jt6bXvyeZ0J4Uh4NJ16efjdqTFQei/YEqgrwFXWDKyBJPey3W+jg
51gF6737LaJo9ML5cyryOsz+CBm/Dowh4s2YCHKLGokUOGvx8kkK45SCqsCUfmzOkiGYVsC1I+ZT
Gan/qmhDbUk0GrGL2nS+xozl44zCH3AoaygGgl3jALKsZblq+apaQcg7G4t/chB+TwKsGI3Txo13
5Je3QmOnjsM0vLQjThIlsg94hBHBwtXKvfiGClW+vLnN+rfJu3K/roEgjoTVn03u0Q+XLQtIfAh5
+Lkd/l2QHB50BvMDHurWPA5QrDhhGQyoYfTYvId8hYhT3KyzMM+V19V5Mz2dCvW2CIkXosZTXH8Z
6M25CiCIJcCmQqGOMC3oamyTGoAUCD7bI/WxfGzKbN9HIpabL+YhKKZHKI5J9NKGBy//soMuoAvq
gfmFGHxDQwUynk0O5qaRl149NA/ElhWG67y7zz5WAZOS/hds2SK3KT41BBoFFwz43Nx7LbJxwWnd
/MJIoTHLeV7STRG/DMd1hq27EynxJjAduJ61t7L+Nnfyd9yEUy9MtXpD0CYUyo11r9iTdfcLj5S8
YjLhc2oShodg2E29FN4yBMj+y86n0tqw3jGR3kHWGMe1ibuaPG5VnWMtx17Q3FoMkCIIcGWWwSe7
JpBfVp6npSMcD7NlpwTrBLtFmpy3k7WSaNr2n4zY0HqynWZyDRq3m0QONJ4DbvRdrnlG+FKIHhRg
vOYJZs63wZsIx3+97USiL0zsEtuWbTe6boOm4yDdcgl9SFnIM2g+3IERjEubmIrszb6os1qDsc8K
l39x3MOLsZqQG3BOLBKQo97dsuLRx6+NZr2mc1GMj1OFv2E6EWU8KedX4qZH6tnzaMgbkCnbx58n
cqgHSHsj9aqC9UVmjHS2KhXp+GP0Kn4AGOaMZPe85PWIkESfgBpr6Enl9deV8odNuI5axR0cQfdA
oIue44UOcEjf/cpGAhBg+W0JV82jBqGTLTmuxJtC2AKF8OKEUyleOXd1xXn5NMzoApeLszSIhMnQ
XUQ8JkDnWgFWsRoYCh3FFfz0drWZPJlqTHjNcDcWN8ga1r/jBC+eDfemdcBQXn0yDHWOGoSTlzPd
C638Lpnqhk7hGcaZc0MytuaG4XHh815VElZ4xjF/Gakf8MqKvX4F9p88LWw4WF+33JazAlMilOfb
/y4gOeXin/oDACNNOXrCjj32QwRFMaeyPUfbThlHuGdBD2wPtlx1XDVb8CidykAC0ro9gO8NwSE6
zNxCP+XfEthDzcOM/VMZfzlqzPJfInV8Q7bcejrPCx58jxAl0hrzLYcchTSsTdQvl+0WAkin88bt
rTs13Smp5B+ZeV+MQWZAXCyGN7B2/qlyTM9CPB70tNi2xer637Msn93hvfWoiohD5+WTUMSwKL7+
NyoxbNWX6wTpQywPZcRosZFUm9i+9m9O8LJ4sKhyKmTQG3zpEq1muxsFDlHGBnDzXQCbG2nVRZ3m
/jyTXizdoLjRpsp1rwi2S6RXZX7iDvn4GYLuewwoQa/us2lPYcbl0i0vB+bQPh7ouJGc0V+ms8pz
lOvwZQB0nPYQRUz2uYG606rBjBlT0ha4OonLkdXNRUD9xlL6m2DzbFmd8PV6l753MLe/A10dkUB3
fGvkamtGYzFgysp2uwTMPD7fInnc4hZnyae/KlPl1Lx4btJhnWmXYPCjmkCrg5lpJNAVm7PpcUkU
RoOHTLwPxWtoBC7DZ18K2DZ2NNvvQmLYbAMetxs4MTtijcQjOHb5lYvshr0rr8RI1W0TIYJqo1pV
1C8zcbrdRuknIa0fgTBbUY3ExMxsZJ5n4MDzV8FaHJ7TBceVdy0IjE00Ah0aTIzsTsGBlOEaR3FE
zZXd38soCZ+cOCVBlz2t8lNmpbKOph+dCyuNTIS8O8QlFF26OHsbXH7/BiMYySH3yNXAwjM8zRHF
pUqC6NpO2FskkgTRD9+/+3lsH4u8K0qUIkjlOYy5SjASR7VWLcY8vwZwO26ISvFp2vjlbVs7rENI
ZLwdBhT5SS2m2xzuG7fphmG9B3HvTj9NLmy2zgBXc3SIAL0mOzoOrLyG+nSfec53/q0phqcrUQx8
V4VQxMlhIEQlN6wHlzNKC37xYwvmeWNnqtmB5fx5scph2xihmkWrYsKIUoG6T02bD6d3rQgunWr8
VNRa42b/MuppKH8eIkq86Z2UFERL63fvkLXIIRVflr6n8cZoACb1q871shb//iIeC+ngBZLbCF8q
O50SeM2beccQpGlR7BX+G0d3M+ifJQfWwWzSFsc7gbRadJirZiq+nn1Hu8bSw2ManaZzjhRJd3Q2
+iOVkiL/GIGNZQ2bOpVhlD7voxQ8HVR7DWDS0km+nCyJISx4IWe8VWDaqKA8Fj7LY1KyJjcOC7f4
nDgSwqbAt/kCFN39VCRc8OWFoS8Zjp+ch4mdLR5tRIVSC5KQyB5/xxSrkzoDB3VBRJ/8LcLLDhQD
LQ5LrTBw9r5Y3R3f/TGAOxL/YLKcJnmWsEaaPcJb/frg8s3ojWhOCwjsbux9N7tfSjW+36uGLQcX
bN01zASmgU0K/sZ++6cRUhA0FFL2lKxvQY3JbNo0Z2p34UHjUl12FV8Ssl7xXthrryYotjy9JA3h
4mgr+qmqX8YI5P88JbFc6+t00489uPlwgMKDJiJNBvfwylujSurtyccuhEgzK5Hq1ePYyjRVMlH3
oL5vPwMyu3xI/CQjjrtmJVxhI3vxJgmDqCXbOzKLgYptLSpSjV6OP8WLKK0yxvw7bVR+VC+Zd/rR
2b6IY2MXp0lpGgxqt7vBj+Z1t33Nxq786ZTXT4qdhLxwrB60nTnpqSre87OI7Bd6xQgxepOyJ06y
rcBBwQdHG99GiSKqkWyNzu9TMc1DEVsCEca1/xOpv7lplkdALfLMStH2ZdIeSsqH3vvM4Z2bRd2N
sPonzFoND8/MHt5ShW9FNVCjdAX//ZGLslvDAisquCtwPllpZ3LbFp5gLCo2FKdHXS5MnweLR2OG
Gd2rsOLsdbMjl5iSvR/h/oTNG7sGtlgjeGwU12j1DQAbuCCX82MM1+f2g9eW41QXB6mgz1Pkn5kE
PYgfZC3thqDx/L8CWYWLdMKJG/oJ6MekfIKyrizRmq4qnDNxN/4DgFGmJl9zcoSPgAFQyi2QHawK
x/x0tqRvH0w+AfUroGZLtjqNNF8Nv1y2RCVXtjFymXJtn/gz5UBrrq/IvLxV4pzuSPUKGMntA9iA
D9FsX1T4fPVqo/d4n3SBJ29qM7ZoLXLD9wE63wZ7wAtOm3nMwfXM/2actG0jk8ovyCpzEvsfhSaA
0vGly2t7yXbLTp9vCTN85+fx54pqTpiSq9qL8XKMZJDrZWyOzr6HH+aHbvP2kfh55ZVbshPVHMpw
9zMxX0nyvxozNWbEcbZRt2BPeu+CHLB902HsKDh+K2owb8rk8EWz/71m4Zdbw7wLoY/Ps0Qy4x/3
FFH5Lnwpxj2bVSNaBdU7MAV2bOdNeMQkq04ebC7zqi5RBlOoVRZslPikz9d4jOxsBvcbCuOJusCl
UZrp6vU83napc9cUyek+xbFcATJFSk4XXtM9Wvv4F9tkUy+atUAwQF5sMRMd+7aVjCuSwUnw7YzR
eyrow54F/1XGjRiaL3FTY46L7+idNvysts3WejcYTK0XDLup7lkO2tYfDdxc/xaPRjpAJtXc0LmO
50gB7de13NRpzs/qFf/2ch+3cperuvWgzJQ06xAaBnGRUYTqjtAvYhJjEJV8mALotIfCNeqLV/tw
obOdvVNg2jbeyoVbxRLB/K9G+TRD/QD5+APgePjddZ0/RUSHKaumaQm2107InAXwv4DJGY3piqIE
iG050dY83XAHmmDB2SaxYYnloDc0XgHDe+53rD//G36mFeNGGRcxKPC2aIYSjLHv2qNuQTaJ2wO4
tNk1BpmhR5PIC/dQfslnG3wgvD+JoDBxrzJujojEGkzKPMwTUtqCZnETDnHEbpuooc4EPvqB++Cs
Vlg/0jOuC0xhi2odtPq4ElibM4iizjZH/PA+EyBoRIoNf+32FJO+xMUsOmnLmn6f0pY4mU9bivdq
ZZ6Gj28JHLoDcrIBgo5noetCu3+WIPD4bU9M3u3wIc3gPzOaZNTEbWunJJJL3AwZD8QKrdAFGRzZ
3QxJVVtMZPkJpRSVtWIlvycdSyk8z/b1+z+pzjCgPbhSOP35GNilWTgVgOzqEM4z7pmnfgm0NTbp
STr7PX+HrqPzGjrxLlNfe5+quj7GQ/r9ZfwKMu0A66bVobtrh3dig2M+PHzhfibpk0H0PUa4UNMT
Uj8b6morqEAA+CAOppvqU3Zf6nVjC/In9E6aLT52IukXj2mxBB/Q/IuDyYXOHsSoSjxQU4KaB+VG
a7Q7CG7OKinMS6DdN3NXLsTybpW6udyOe5vNgBnTN7m03NsrUUv3ZR6UA7N4BAJwXMNWtfvkmTDA
j4xObyyHEy+ukFRcCKWSAq30wj+G6EiRU7as8DWFSoyKXBq+27MMR9E0HB4PKRqXeHuOlnpXkj+O
Rgg3QnjoFrEqmL42kVuyz/6JkotaUo5JqjRFxfTmyVvYHFGm/M/i7a8k0o9ps0/SI/OFEXK6Mzfk
zLNnIaI/aXq38HQgd5sseW3/1LKcUJeUGTo0NikXweEsgSPXFohS44PjDhjfKOs+1uCdLr25oDDr
m6mt4+Mazu8zsH3KvCIMxafjAzevaMg6ooPIQQxGsqYOHNWr8/67BEKvCYuyKgZQAcdYmB+qLRFe
0mG9xNcbwqo11GikyNx/29O0i+OUDpjh0Fe7uuAKWSrqyDjJXOxf4ZtNTUuIKhq613Cj5BKlJwMr
8GAeNSV+wLaEV2Xeed/s5b7ur5WZ2LNxZYHZSIN8uCji+T6ugI46JuIUS+ijQOdZbsH94umxuVhW
ftbL8+ZTKBPVoN3WEiTconBv/s1nEJ8/ryTtnsyWZ7ecJK4II3Hj6wS1A2VvIh3qPmeRoF9khbZF
OCt97FvyHvqNXUl2qFXoSLgIbO5pEmsjhAwEzGXJPgsecVQ44miS7jDf8+DYTgHMcilikbaQnHvL
oAguyd29lGVBUF2pkQURsOOPOwGU9DJRzFdlDMYWpp8GwO5jG8IXwr3vDUDax5hp/eOT1K0pFaq6
PK5LY0NiQD7ujoEgUUl+RdO0ncr8GIfXI4cqguKjoMgOX2hnzYajnoRv1rJMoOUvBXK7rmX0m/vw
LW5fskRJHJSahZrJOnmfXWz8Snm6IsX0nvAUOqIBaZlsnwqKkcn2kCDibZhmFwigR7/N9dwD7m/i
dYz/ga8a6ZCHZNl50NTfDntnVg2F1uNcLW544VtK5WNU6rDYkgVwKXYAFq1h+/DFf1fUG+QnP7sq
3YLwIOY84kwkFpFo9sxwS7FVHBDP+iO4LL4krDLxPUUAI5HFVl7gaRMYMMwc7WOy7DSqjiMvQg9v
1TwMQ2cLolvb6pGc0hpAVtmeZuHpKFIk/xi2a5jcU6QAATht8fx5gQMuZVeoii9w/up0gzG8i7gH
OQOebwonaQiQF3l9SLYpK0vYmnI4PGsnKUwUSNzCoszt16fwS7hFrTd392my0dUf/h9Sok5p52Lt
9zRB/DMneIrtCPVNlFUI/c0SjcXVvkBP9IbUjVxGBcvyaWs/xFd1RIsmkB3Iq5ofOHvOv9ss9/YJ
U5rj3lv+r5iyTYUiyy6YoNlkJa/NIZbXq+YLwHgwV8Vmf0iucZF1bS7YcLD9fsxL7vurwx1nXgmq
LfvRmaSzJQVXpcnLHAm3YUGvIsHfBmB4f83A1gGhjdH6jJkVqr+4GU7O2QBSQXrdusSxQwTy9Fpz
ilFzFCQxbZw+AxoYOpjwB89Ex9n/TEfkkolGZF9qy6MnFJa3iFAu7oNy7Ui/VIIYm+xR8L9qAfYo
yDCk3T0r+bG1fzuohyfTKPEbrXOixKpYK5jAK0tpksWtMb5XzajU2K0x0jjURw7aK5zyKhzjRpGf
pOJiR04mo++sv9bw0lkcHvv/RMe5gaCz0DB9XY1sx5stSzKNi5O43DRXK19IrmVnzcuHMnXFwwJo
iXrzdLGLNX4YQhpNH6pnSPvKiqXbGUyJ9PtNv+pwhDFCQ1zw+IePzuVBKEVHTMQLNINAFrGK8iO2
aKxLsdMCTOFjNL/KX1YE0Bj20FuaXbqzm+YbX4zGPs7anAjkwMB/arIcjC3T99wrWpb/7ECVzNVg
pfnMos/owBqqyYHdKNPvrnJfFGP1feFMxnf1Y/3To0ksrakyMKQJwhYpnz9rn95REl48EFo4onK8
9nNFObZjwnzpOPArrMWhxSrSCpzPhkILkFu2r6luZRwnrpDS53jPOHi4jle3OHuGIrrUUn7U5PYz
FMXUn23RmWP+9bL/8cVDdezRkM2EKNdUDIODWYo6dPnCpFMVT4xZVSnngK/XiTkrWwkdkik86FUk
8eTJ+FYrTJN27utK+pSf3egXocyM13JFELmaJygkqbV/6Ihxk7148if2R4m5ayCzHPInSCXUJtAV
IuSgIjXiRR7SSHTNOSlqQ+K4IJQOcBoaxlwe0HjxIMVvDUzoMuqDYzd6Kxj+HOvdw5w3YO1tq/gP
wS8y1IBlGDcI+YDinXzLUJdn6UFWEMYaDdBMj6SqMu1KkzqMsrDtBL/xBY3lt+s/0/YSditfoVFE
wvxT/HsGSzeAmM+/m3+RtEZZGrYU2B+UROOcvcchSV1Q2PEjJ0OuQJAYkQxADnviv86S7Kjp860p
YmnOLtEvuc8o08rcQgjBUSUuORy9KL5zW789T+vwK2X1gpjjD9pJIHCZN98keF8vxFQ5jZZJdl7I
+tY81Cpq8N5My5xmp5IR5wEm7u+4P95nH3YBy5018k/uDI+ytka6eEg/lSsPdopjCp+IX/pwRTU0
PvPLsTAiyXW6Ea7UaqEuJSxM6OzUFn3oYbhcVHi4YuxXbib+il6h6bOk89iE2p7s1jdu8MrBMagg
SQO1hKXBTHD0k/OQpVUYyIPCAajCmF+4LJsLRGMNAmhWNAECvyzmZtPOh5nfd6vlTfjDYHwHeFr6
w4FOKjUKrnny1Gj1kwj9izGopPlF407aKCE4cA2v1LmnVINkmBtxZDPrwyiOSHVvTIYg9L/Tze1l
JaUEwFTn/kPsqKSNNGYNTqmQqH5iuvDldY7fsWL4zao9yDWQgqPx92kE0S1bcUNtkYbCoaymF9BI
+MjwTcjV99dv0zBvdoCG3PvTd5CuVo1xGBbBUhdMmlnSApuE1/P9HSd5/mxJK5Y7omoOw8j2j7hh
DN+ecyiEUNgsgBv3TiBkGWcRr7Qt0hPT5Rv/xiErnnssKMYNPx+0Fc8/NEv44rgOkV2QqqcQTxfp
L+OAzn3QEwgzrLjtCyhhnnI0Pxd9eZCJYzCz7nZUGzvNYp1x6Ggwxt4G4Mb3mCfVXxEz7/fdQIUi
Q7h/9VuG0I6kHACODmCUBr7pAKRktS7J0d3Z6exAjx7QUWzmXDIIiQctFEjGEeD61XSM9s5yPx98
8nA6D444g6CW6z2WtxpjZ/Z+6zo5YmJEVq1+KqBS08pq87BDrH+9Vr4MfEwjv9Ru9eJvfBQYNaJ9
woT4Onb7ekCroU8rESY5yUyXxr2srJWhQMsix/tNf3kHFVPTTnvLpe3qdT+BaRrudnFL8Ass070i
yqKjEdp3+61cc80da2C+c7yNawNt81+EjS5drYiX2h4hPVteFxwVY5aBVmMZy+l/MB3hrsKyllEJ
iZ90VER0PbCi/8IrE7DhSuQezECdGMSGA9RQha76CblM9fX1mgomEgDbWDuLoWNVRNtzS/oBCFdg
PgmboKXfAXIMwdF5xP/RmvDunb2m0KGpuX4KY790c4OU9FGcD+oK50Rd7d/SycQq8ELd4pEB8sU5
HqkBiOOMYl+5eUgwMF/upxfOJQwzMUWY5NsCs3yHN+GfX4Cd/zs2BZMIwgY5pjXMMtHcMzZSvv3m
BxRDOtNlo6eOylkm57AdY0hKhXLVj0VFFwClBWeQ1HuckrpJ/tKeZMlhlhcCbqMlOOCDGQcNDF59
cxi4+H2a64Z90BbN8pOQP6gQxCB+A5MUVHcRAy0DvHlOJcRpkT+KV9QkTid3/npCIB3Ubqlz2piY
4jsPV3U9hgO2TRYWQL+0kHc4SFVz7OISJczq4fNKJRqYPYvzjf0Sx687JLz6lM9Nrbrvgt6+9krd
+zvjrGIIUCeL9+OFUV+eSw3Y6kLxRT1Z1iSUgPYtCTxsti8UOw/pd5BME1MJXhyWuNQYod4Vk4Ca
Dn6NoEk2tNmcncV8tkBWUs+RhHAx0ukzAvISFj08ur4Piz2x2+U9N+ntqdkuRuDQ1IguzgEum6mG
SjJ+z5UUx5krgT+v1plYVTOpDiH8jX4+ubIAb+1lYWLEMB6FaDqJxK5qX7DIgVcSJTRS8nfHBE1K
XE7oem1F3L6cW4mgImBoyTM7kjNgoNKRtEbVbvGzx+g0EQNygHjPzoxdjkai4vygne/xdjNMu25P
hOVPyzH8scsILelSFTb0BoSbzsilIOTzSMWQDgukg9uW3E4+LdavNKmEv8R3XaGcUGd3cIMOt0Mg
QA8L0CMDu39fiWhidFtKHFc0z/JRZl/1vU5avpb2sgmbiIYP4Z+JrqwGwXbMMMSDMbenmuIY1Egl
mzc7h0upn7PGKGwMtTn7XzuF4Bp0DPFR77oyEKHU/ZvoofME7Eih++TdIhFV2rsKoLuRiUqNX5tT
EAiI8sOUBYGvdVg3CmU2n+oB/Mqe5mXwX4lB3lCYBvd9d8CyM9a61a9bLq2rjoDEn1n/oU3DSusp
r+bG2d7ErxcTr8gMz9ua52BR3vnA9xfXmNVPw4eVXSShuDB1SfRju1UrTcNUEGO0Hvf0vKGmlVAd
mhkMNwUsDq3nNr1WW0/LNKHyLVZwp7Vn3J6C6yEXen9uEseIZtlF4v5lMXl0Nsv6jJy5ZvBocZnl
zfMNpz8+aew6atThWYo5TdpJP92/KP68bA2dJGiuPB2H7gJA3AnRzGtZnqwUQS4WYQZlYzvQy0RR
NgDdtz8NHBcJqCvTlGFFFvoKTKRNnaLeoH91PwKIcxgMmFaBovPkqUop9I9SfVUTE7BxHjJR0rqg
OWQBuEHp5Ju9940xqTd0XqEdaPBokJ8QVwTKMDlazz1aSbkrh+MoKlaGkjyUhhGyghFDRNu/YW6b
rtCAxzMqBbs3JOM0C16FCU9yoobOcP+QDMtZRHjIq/EGOE6aGZYQ+VjxGw553wiznze3GHdqpE7i
DiVC6mtEyOv++z8sdcH9aYF4hBmKvssmZRnIjpp8fi0fnfc47kI2UU0yZdCdE0Rcs5wDV68mY9Ax
if53VU50dzFbz/ijMdM28h1/Zav2RjksOD7+BDfq4ds5Pl6yDbBGmJyVrrIEdOuIK032MqxMUTT2
Ec5D+QDDKSHYX89yPyfZbrJuqxp/1hqlg0o/4pgEACpeMLP24PDZBoiixQmW3apn8sZdy1o9F64s
d+hbmOAQMJBQj6scwAuD5ohcLedZAS9oU1LgBgmOfzaxkTAkEoGGxK1omZyHh6MC4lcEH6yFjfnz
fP4+OGEnDQtiuPUrwRICq8oQb9pn5arWJeffkiOTKT+ITwL2IFXPM/xm0QDidRjqmcuYWd03x1vu
I/nbn2Z9FqcnsYYVefUtmABILi+HQ5fOcun8EuPH1ZDed3nIfL8UZJ+ugRXjtLTxFsMIje/A3LQD
Bh5SN/nHGTg5OzUQyAhWhztUtNSUrY0Z5fvJPx7141/9BROvl3L0Zznbw77j6D0M/Cc5qLsXMnNl
zZVGC80ef8RUEXBSUfvi3poPnjIzOEMgjRWGPEx1kAChEDEdiB85TgWrzCW9z6eOEQs1qq966mHu
YLkSWJIaJL8mWICJG4ohXi8QSuZTA0sp6iz96dyLlC2vFRLxWGmBE4fD5WH8yAv8X18O0cxSex0a
DgaxNjcQxEPmvJ+Hp6PWWhJ7qPuB8Wro7FyIgfFJd/OrkqXGbIb06sBeE0rAuimfxF8ahp36fd65
AHb00WoyyqfZlLQBrTjtIrgbAhBZqjJUNXrihrrqhh2sKhlfhCtOOLdKSiU97lL0Br4EzxTVOfD/
Y5Sf67VrdNXHzUp4ltGzByIG0YfnGRwnsL8w/rY5VEYNf6KXlPZ2o9ki5FesrVNSUNf2Lcio/FRe
IAYVQnPECZ6wZvaQyfcXDnJjH2dlHQu/oMhWMFamCgpmzvnFD6QKKC9MeLxdBJvFIeR1+UtPKmS7
I1CYO9d8j3S7XKgd/Z13gbJd+GKsk8JGAx03+USgzb0E0ivMtEaN9dfSh+cGfZsrI9CN9SNYNIwU
jxTHPvkycLedH8MOee2Nsr6Zxdz8e73fWqrmFcR7mNAD5h4/l/c4b7YVyTk6bfmSaCGA9+g1x+Nf
pc7gU+8Lxu3N/yKgwb4LZLxIOAmSHmTPfToYb/vIa3n5XBJCLHeQSgNz6EX+sEB/AWvgC+/VUY/y
RNgck1M9WNHs3ljRr5KfN5IHFVmsqQeEE6I2BlHzpr4KITQXBAjeD97kVsG1VKVVNV+ljqKFMQiF
+3h8K+DO9b7YvuDNLSQ31X8hs3OmlvMgwpofjWxZC1YEmsdiaSd9KYX2gdulx/w2fVhbShfH1LTn
d3e15noZjn6ZNJdmD4Hj41HR6fSVAQt9fMwjPdUOvLroF7jOTE9MvlBybF+z3gw08MDVvGbv+ZrP
vXcFuo8buCgk/fpSb5jwagN5f/qnVt6H2f3Azv00TrEHMNRp/V5YyIRx85CVrmJuh3N3oMKFKxPv
+/zhLODeYk/P315BYRHI/ljTsXMPBUT0InvrDgM4Hhjn6o86dn0HpFw4grLPs4JOZxtwi0NUvbs6
mam7yFtfak/w7XmB/uNlZcTx4bf/zVp9SgD1o8TMgxejzKt7fH1XyHQ6sOqPWXCe8u69ru+FGrCH
R3Si8JtFCn74tIDsA9bPxymeBphbSCSR4sgi2Bz0nlTaqT2TEsMGpllO09GhGLWkCpw+X6TnYVAG
gGni7Ny/HwOV+ftTX5+0qYtq8GO+A5zfkuP4GAsPWWuQAeNIcWjh3JxiUvqzau/v27x65eVJQHaw
f/QKTSqupSoSloswamtDRjaaJHzg331qThyQ4VzRSbR/wS5cavmRtooSnvUUxlgG9RtdGOagSXZ8
RTYiW5O3tFXs6tMZv3xSZCOAe64o80ssmYqvNrrSSttnKn2vBw9uNNat2jTq0XD7UYvC59B+A3bw
G+q62j7SP/MhWA4RdQ+W3oXTmpiIY8gi+8ytKrff3Y2o1fsMmEwwf9eatD9EvtCM0Fv0vaBb09bW
FyBej0DN3MGH0NmWn4hvifc3OPAEyS9oedOkhbkHod/FmSVWeGxjymdz75982I1G114yIjjdcI8r
LhqqXhmop3jwZZ9sJMmuTccDQAUKDO6MfNwhfpS7jHQlYy0XGPZPMDYghpA5uuen+l3ptZQrWG6j
B1mJAW0DEe2QgokrnKSG8qU6KD7wiJxWOhR2Dpm7JDWERzrRn3YrG5fA+q/VCYlT7H+xCM8x3Lam
i5qcqc7D8LS7U+1FcZZSrtmvu4bcH9/0VPvLwjczKRqxr+lAuejck2q5o5l+qRg6VpoYjioLraVs
wWA4H/UEMJ4WKUdMbhkEynnwpsuggVLIU97a3BSUB6SgsAFqcZIlbq+mUOR2ws0DqfACMXl4gE0M
I9EIeLb0kjpaFs6yzn1i5qju73bo1eHC9xjV6QXRv2V0qUExVOi3rxG9gWihR5bL7y3cWXLxzZZ8
iQOQxmTqMK6ZQnrDIpifjsV11mm0tSxs8mcIui45OJJ2PbXd62fpO9THi9KYu91nq9TZLWPE4S7I
FC8OlVFI1YY+BXDRgAh9Q7/vlyXq7S43g9lqjBkwm9ob/PbmQh/Bk45wc+ZMaeNAvX2MVM5g1JDy
gd4P6LMZwN7CEOYJDolzY1eonxiqtXFAXrcf7Sp2o6NXXkkn4uy0D9JmrPUbL83ifeBe04FqHx1a
yD3L2sMg/xXQJwNZduvih3epGI5mxPv10Bj7LSuHT5LNjG2bVnuntQjTH/249+MsUxDKHJmwiiII
g6bS47nxoIopx6mZ9dDFoBigcdAeylYM2wZFTQ/dgKfwwOdu72t9Nniea2+m26vfb259IwUwUUmO
9VMu2//1/wrlm/HiB9HDer9hth8tSaXN1J+elyLZEurUz475TryjP3xIL/oAPLxw8w1Ygq8/HMvY
5t7u3ujcvXm+J1vVrzglGq1o76lpaXmAnfJoApX0In7vuu6SIrP2fwCvk+KxjfZgztAq8mMnUDU5
QyQA0PWZqWyEh0BCaucbYn/OBEu2pQSoQ4eWUDgu0wH2TXPVIGYTQfXX7OWv2NWDl028LD27Wav3
RzPDvrRSbeghp3cK515Xr340DhxkbzgVnBBfIRr9P2VhhU+3Rv4OXW67zb/dBtuxfN2z3/3dT5FJ
ePGPN1W9nf7s57ojaurs2EUvEv8ecjjw3CVvVVvDBbYzWkpxOR2iZ4wOge2w2VVHAvEnA4SKkaq5
0ChrgF3YRlv5GZzBvsZ19cQPtmS1aof962bj9rocJiB1cMKuYOyd1qrM/HiowCl8iDlCJLKeyoOM
bTW+t/Qh4yPPaA8DqfWdz6WWBPcdSMr0m3qU6S6EBaBxgYtVAWISIfEjiBp7mhNSKt7PboyIq+1k
iGXmbD3RD6GExlkRyvNRoqFDGPBcO+RLdoYB5c21V8qD+YT4IeWEctp7rEmRdtFaG9c2kC70OI34
j8AVUPPuiAcFr4vwYDDiMafZGyYzlbfanpUUcAQNCN2ZusRTCc7QDHJhmP1/2kfS6qV14UL6RhLW
8utrJwnVg8zBiEgoiqHxJl0elNbmRONoHWdTsILzGhCsl0H/7cqUBWQPdO3YQpjqdVdAiNzt20sK
t6suhULRL8IU9eFOtN+mkGZ340JnBfUHujCb08NT2yP7CHVbKq1XBjEe9rr7CBv8C7xOPlKF+jOC
F4KwCubFdSLvZyqisRqCoyJkOA2veYFBI+cgC4oUJd7wggeKqAogLapPN80tobyq6okUDLr52BM/
7u4vH8d3ObOufoEkovvjpXgMHKzJVfvn17VzrzazjNk3nSxerlksclaYk05WQ81o1wKmkHajmeiT
0q80m0k6BKRf+yf/SvypzGIsjhDRWJAFkj9gVmeO/VaDErNkxJvKfwJYSUZBX6cp0vHgb0TdaiKD
Ss2oOjQ7/59WlpVjac4+iVhZVwoR8U6vizNtFfU9BDFZhnn6abu3b7bJuBgz3AiKpRsfRlhlDQWo
zHu5pDVvs88QdYY1lv2yKySO+q8pxQ6B4XUWsAerghXu1wtK6nNXRErBSo99nNbPEjLmNR0SAo3+
D8jgRDHC6GIK1OlNpxFo5Q/3yZfzuP4wMim5+kM/LngQOt4CY8bOQloA2mrO+FkEMT6Ee7xjb7KM
vn2OFFsDN2SZeGX63/Pix1RTONVk14A2XzpuchwBjyhqKPDLG5KdfoaYa/mUGVSfG/q7iOjrWuus
ntV7HX5Hw9JiYV/yn15/942lR0LEJUgyjeaSa6bLi1F+TT7Y2r5wtr9f4+YwsrbZmLezDswO9tqM
i6DP9mO4NRErriT/VFhFZDoQeH492F0fVnXNlbCbj8PBh+2MvuoIdf3Hc3roGFxxY4ZIAgXiyuuy
s8XGYMnqcPJ7OVloIJsM9ag2WeDju1YaFWuYRJkry3WiJOqCS+HmRfRECteW7yD1yHBnxH+cl8Mp
fiYikuVAn9a3/4Z6LRMidXFs8ODIMWzY+s/uPK/12HKQMvPxmYtAOGh4s69ZGfeuNo+vEwaf78Q3
JR++aeGS75JIkA7QizjcA71iaqqCtJpf7azZoiRNc1SRsrcpYnHFYBE7M+ZicPplOhswvZ1U2LaT
2imUabFAmlDiVjTupP7CPqkVenqcXLAaqsXowvIim90nbzAXca8tDTnNVldVXyV1HcieFcR8a5ZE
0znzL6oo4gEaq4excCdQfsorbwhvZB3WS31iOcbL3ZkXnQJieSkyIYOFaDieqKpbNoFEmOXUMbrO
OaHQEa/TVWWAeIBW1TJWa+Tr0kL+KYA93oa51/83E6sB2B3Y5F+afHLwgJ35FmqXkFaGiDznLZac
CT0HbKMvMDrptsX7dE2+X2rE4y2Bjuwibl1yKiepbHfmfWFU5gEB7QT1zT5DLfPST9+/CGFuqksg
D0+yd0v4gLR7sgd6lwKSYv8N0oQYZ7sGWX+gOQKdtKxLS/bjOVkmafXtZ3hAtP4E0ypnmFE/Qimv
v10OLGAoNdsTHvnZu6b3FISNFiaHKh7KgHgUwNDZGymbdnjtP6bmItXSaPfrFA/tcr7KR/yZ/qWh
ErqiE9zmuTsRbFFOjP3RZoEAHQttwtMxS5oD89BYVnchuuU7+0uqnZ2cKWO8UCRXChtuRB/ORebf
M/UHDNSJCdW//D/YHaou0fYLZrbo4C2U4DwY7eAMKgSR6Lw198DIh8DuWuz1JlUt7xEQSiunImMR
IIamHFH+IU6rqsz9r8V+YsEdzpLI4zp/cNHnvq/7JCrID1sV9e+q/F0BcIwrw+U+VwBYNIxdrebL
gIvBAjfNGD5rSLI7gFv/gYKqIzaDASx48fFSzCaQpOgg018i1tXFd7xh8qBqZmL5pMHu6Mb1bEpv
8dvehM+5S75mBISlO3ylFg9hJsYfSwXLj2/Xg9ZSeCA2Sz2ZrZKMe9pt1XWhhFuJjA1WpKNr3oGF
RhqmD24FrbDelA1Edu2+yOq/mGqFrJ8pj1yn3mJIdNZGnnP+KYHQNsPBh09wAmWdWv3Kx/ifEK/2
3X00ec0kLH0uVD3o9Js+kb2mP224s6YPZkkBYhvu+eR0HriQCBS87Qo/aVT+H1SzcgdHl908xV0g
Csax5zQLMAjo0FZ9wrAzkv97p+9O93oj4DMEh5mM1JHD+IViLJQF30ft6zSaXYYzoQphHCXhqyKa
w2laAUeP/M/rLvUnfvPwdi7oGPoKn6QedIgDOcgoimH0muYjGx6VucTg/70s4g5tij9mFi1uRCaD
3fIjbgWwimnfdimfT35Z2dGTJAUh9jaYxrk62qx7o+7uqUIJCC+G3wYndopBSiOwdZ3kdWZhwP82
HuskLhdD41WlynsP3rvpnvIRe3ZotffY6xxWbDJezjnew+IQa4lUinxCUIYGYYwQNPJdfcWDS+t3
vB851HoxiiQ9GqW58Q3YF5b9I3L6h7mMxUSRNeLZZr8L7GM8x75UAzZ+k6qG1mYUM0grS1qgIdbX
sg3aquATDwmkxY4pHyAyw3pmBDYngHkIRXZu65C011DFUVwqSRlIwhVmlnYpQjFy8fCOf5gG8/Ri
ndJAwqu8bComUB9l4mvmImPAw6FykGOzl/1B/Gpz8m68yvhHS6LB9/lTQ0Fq/3eAexEg3pdLQj28
H20dPvG2emA4m7lOvMsucy91JR1nuGtgA80fLU7JbUNjKlQ5mAKmGWjMkhXtFWd22L5BblBBvb62
GrUgjrZ5M9dIRZlw8aU27cxdwjAcaVrCE8+RJ70IOZBeQXF3ltiKYe59uIeMMGGiM0l3mfgjB49N
TAB1UOzE0CV17Fui52vgNyBtxATDE7NNtoxiMN8bmhH2OQt90JRvyJ5AsdI7Hr88/cFLQxLtzHo5
be2xvATPoCW+2fNMyR+QYMoYngOFfSq1BrKKlTmQe+dLMLOhDv0WYAxW3299cV1Ve2Qy3BLRW577
XiEYtz0Fx2aOn5rGwYqtO26V2abms5TgBY5HDgFv/tHgtbsTRvh8QizqrM3GuOA0Qc9WoDY+EWQl
vc4qeSvsWGOqeGWxvq4492nO0oWRKercMGJi9FA/+pedFi655+b33U61EUXxnhxcBcTo1B9lfr+k
Z8N0kyzmZQvi23Vfrd+PuP2A6Kh1MjVrwfw5IPq/g43MP67d97tBs63SJLzk3yOphjzhJA9WH9SI
TUQsLs95pplyltAuZVeGf0sDj7OSnKzKQ6PnkjfZc6UT7M5FL5wgiR4m3Lvw/ymT3JNrAyO9vEr8
bV3Hx6esJOf+Cj4Or6IQyCX7iCLHUf7e5CcFnpLt5YdDTb520Ko0kPuGWn1uVlW3RN3eSiQ6phjW
6RDrYo9xFYZfuD+Yi+dTwA2j7d/mfmChr7WYsWuqLPHAqSYiSI/56nmNXa4/27wpxBUY0KKxQGNo
ko2cXaUFzTceV85LUugogBeWt6bM2AVgGQUGsDPv7GigEzYVy6Z2Epi8FsA+smdVCqmczPzLDfpQ
6nm/DpkxDKpdVsVk9mkEoQnFF8lOdGdaHs+sKeYpmk/mAdxWp6jFdyu2BNjgNayMSSc6MpBqe+dA
qkS2WjW7SveyzvDODnQy6kVR5GDpxx78gDNHNvXl0kLxOJj7nXWsBrn2z96e96UVw8UVYVl0O/eK
WrTkEhpfo7RR3lPgARRhuZL2GP/Ugq7hPR8Z3DrnmWJiPJ7cN34KsZdT/1mHHOOEbAaUcPknA+i7
YtZ1/YTsqurG+zDklboRWqRoFrtfQuGFzaTAisCOquhbv9ScwWMLNJwQhtCR4p/EBzmMW/JcDmm8
kjFBYZ7iDcC6TnW59+OXLRu5yhnfDgqfppRBNaZvO/Hx4Uz2j6YCUpz/K/Iz9rvxtDEprk9GOigS
oFjcdh3cwNRYcoA5KlHnJeLXuiUmFPcQRRItX1E0Yn2wpLeDA0DV/DpMm8ufc1W6SYjC4PoHCyam
LIytxsEU7OqMjmyp804+XiQQsglg01SuxcMGAKFHgqx6GsSvArrk8LTCigKvnfDFdwVw0tKYMHN5
3g7ytT93LBhQM1ZgUUEbCPjv3WEWOLbgRS6OSTrnEUbD0TfQOICQPQhG7LyrWRbMhcIkb+g6jQx0
6oEKFXOClsqM/lM81xgEtPkMe2oxpZJ8V/pW9vgOG4yiJgFIjeBm7OGDQiv9F1++ekl1cMHc7Jkc
2eq6HZq+LJ/tBiyX1/bycXI/66WOFNXyHY7z+PUTO9koicCYAJzigcolgXasarSg7UsojMSpd7rw
50yAx9FY0m4vBqe8CzxIsOTUJc/cuSkqJAeTcWKj+cd466nn3+Z1MKGU0QuaSk1l5lPWChgzn/nd
I3lLKomw2GY97M4Fd0shECodjMjkI1Ti6a9oj51lFRhyn+NszHk81tYT+4/p2pYwbN0hqH+GPYkR
nw9aeUPBCtFRRQuzG31HZOCZqGOe/yuva6oqUx5JFLLru/StiFb+sdCdArQy8WHYpbhcjR8RSo1s
rRcGj97YyuMgKVbTo2hcg2yKXghnNEfARj22JcjdrI/3KuAVIGn/3LzT1V6Qii3uyD8rvWIxrXVE
bWRpq9c3GmzugUdAWWz+ypNfn2ZsFV+NKv7XMbdxHIKjNaqoRUbNEAHTHPoaHvscqA/yA559A0kP
Kg+ZrCgCxDJjcp+Uift0k0cSJOZIIo8fFnIHk/NmL9qOT/8Yh49+sn073WFSy8o6h6O43GYky2Gv
8WbJmYZ9SahcluLITt9EY2uLvPOY9DmRqj4TJFK8eNpU/NHuzEFH8FEWZkZa5VY3OD8MCYnnBxJa
fLxMchMclQLsA0DX2+nJ0P41OlRc6uQIEMF/oMigqvGD/3qPncXvdUUfh9+cTTMFIwmwRJI2OKY8
NIu66HjrlNJ2OSBOfyklZjBznXNZwgd74tib7MssHjqtuWtyFlt1lgDbyFbKirBr6rz0j9lyp0zB
bhWwHtkjziHHmulTjsXwvDrbg/2JC4qcU9htpcPmu5xfWYbfBL5gU1D0YyShDXV4FDgLxAm52XtC
ATQCzbVV47bS/8aMVP5aOjUOGR/MElwoft9YGO3Bbq2m2kgApV1HGISg7wwAsHM0/swFYf3/dJnX
2ftt71lCIPTKKEUKD2S7hxBK5B27vewoMKtyvz+qNoFCVXyKQh9+o9gmw6SESC7JaqFu2vQFA4XO
pUogvkf6FwGH+9Hn3H1Qatfk86aPhxlGzrbij/1ddQ9PR6HLNKcI9m/DWlmpUz1orWHpxhEJwyil
7lAsbUqq74+0xy9CeOlElotxHF5nN37jUbqFWeNbHGqBgojxaLz44z/zbv2g1OId544E0w1g9rIh
k+08zaRyyz83QB+2HHSKiLZmGCHMxqp4uSHqzTyJio8V6jjeS+MewVeg5/3zei0VHZO9HDg8peKg
ovPAijDMT9TEjWiN+sA+Kr8oRYEi4Jx0dP217PqQHUKKTMDuVEUg0Lk2bvH7x9mjSnOFojnP4LVE
U2cQBQaQPzsOoy/FbeZf+Hk55k4M05En776o4tXodtiedcitZQiDdBUXj3iFfbjsuOY8XGr4WwWV
/bZ3lLQucHP/wb6u1nOEDZYB8uOBHeb+9DTSKn0o7VfMju5Vgr69yylbB7lAkbKigfYKTaB9PcKE
POXYA3YE4NTNFvfSsMzjA9AFJwoT/MlAjergIUbqUDKWJBPE9jgBOIneLA99/tcpi1WZZlEWTb5x
ixX6bScgyLeMab2QKhHkEYRNMvtI75Agsf/51zw1kFiGvXAiGVQwf+KimiP2ZJ2Tm2Sp5Cm3HP2z
YMEeIfpvz46n/yNTsSSDm5iYjqjdPpxOThSFzv1oR49XjiHRCtA8D4nwtRzauHykPiSzw5YxZb1t
fJ3+OSHON/A9Y2hZlZkboMZSUlC+M9pPMbgSGochwNlybeob0IFqvU7aTDnA9IzaOAfbqYT1d7Do
rIdasWz+syhfSeXyev/7gGqGkiH7KtgsycBzP5hsjkmOb7vjJE3tSncMpoklIhs5aZ0MBaBGDOS6
HNsjDM5QEH2zpn6wnrBFtD8XqSyx7hviVhrRRxrbl2f7/7b1Xg1x8O/Ae59MqfRbbgDdkjFlkoF4
wNOiMXKnAqIRpcNOhENgt4Hv98afGiTAQnVK46XxUbv+AlxRSC3SrD7N56nKJStJR7h1su7cx+SN
Cps9wI5kSv2EWjRZmfwUM/9nJi7Dg/4DcC8fb+hIEdZb2ZquMkaGCb9Cql8oTRwRrW1M8B5c+Umn
CP5BMfaYD2TDPOvlLT5rt8AobQzayTN5C+bGZT9IXbMs1rTw+6Ia08mYJUrbQaQZohzPqxdBC7+q
kKRzrhRFNYYVuCit4I6E616wL+E1UEDqEYgD1grCEAs4at7/VElfrfm7XNYAqI8oEgDJ+3PbZXdV
8k8n1c/uTYJ6BfFLZ3tcmb9P7V6N62p1b7bHYA7Ygn4A6yckw+XiQeWeENpNRT5pvIlOBntT+HsG
o9GQmXCEdZW6IHsVAOcwUMFiFM4nTQl5iQYD0weQLYl6DWDWEACM8swqslkyopFGNTVli2eA5Iui
+t3szma6xUSHkaxTK84Mdov2PZByhGaLQaUEIQp4dlnKwACBGjS62WuEUQngG1l9JVQStYTiJw/f
Ui2NRI6kb9P76P1MA58k7HYtJ/OYrgQo8YXFDBn0QIU7qB5Pt7ynUZbrp8CKXqlRkXbVJ5OtZbCG
SCFEPCclvejv0FYs/yqqgCYqwWtbcS5vbon/Q/7jJYDGYhhQytmJrEWYFibBqcSkuon3CKzlYYkA
nwkqz7i7iEca/WTKfz9tp5qQzoVmTrajD+ZuQ6S3NgI9Ovv8Yo3mAy9eU2aGK5h1KNRnFRSskcgM
lmbrUeTFMc6kprrmc1QLm86vrp+yuwOR7fQQgAdytIy8mNqcjB9ZAPa3/c1xB04DjbfaFj9rvAAm
ZTJ6gEiw67DslIFWusrmanxj4FiS6HQp0hUjOvlIK7voRWWz8x5zhyfwIXYAng4Xabko4jk8GZA7
zEa3EC7pCgUvxqQcULzfZBU0Cd0/zmgFMb26lY6n8sEPrChsnUBtHJOgewIu6DFy3m0cAh0b9DnC
xqm9gDUhN7TySSbbP2EzsAeO1RL3GlLxyH59W2l+OtM1+pwfynwbuEpwnaIxux+gO2ouPp9qgpjN
44vMnnL+DuUEREQPPfCVyChN+1HykfXyU7GexY3UAs8/5Pm3gc0lA+ei3HXk/ssrCwfX8dORIAS7
O9rXFUmb0zVtlgebSubfI1YNjHyNZSc4tYXzm3JjpgzvQPrmkocdV+zneyjiYpHoE8tUDcTgO9jL
/aFyGJRac/p++HL05/ApvbK2CC3Ic8IY8vRmG3KcKYI2oahU+OyBZJN2L5EAG9I0D7SqIKM5glcF
zwTw99IpAbcYJsWdCPO78+M2YrpZPV84fjMkb/ZvHsh3RaiWlk/PhJkCxUNDqN0/cvxOWPP9F2hB
3sjWAeLpUUuo6SdzDCuyCWVMWCnIIWhShWmAVpK/1+oUv6CklbNPh/BuvKkLjHlwN/86l/jwYGlA
giwT5FjxsDFn12+jh1+X2Mt+lr+dtYOqE+GYh5ipK3Q3MKX5ntXKorzsa1tAx+HcK1ABRJNRLSj7
yFjxK1YzDKncTn7wJlU19CR2tHBGMYwEyknz72YMXad5oREttagN33N2cOzBkIyKfCawucIIJIdy
MswdKXke+uwvCwW7b2LuQDF164d8zYC+PZicX2Bh1P2dYrJAnA764b4bfgYJzviXahGFw4uT54Kt
uSiHIlhIxfhdr6ziTmEeHHL7A/eQNw+EQA2BNOQv7+Hs5VkVA2vPxW9b9wAqgQTEYiR9KqTSXX0i
9ALqVrSdFV7V+6AXtmgznB8e3veVlQode0JPdTHSCBywhqO8YB4CsWXNOJuuDG4L8U3BUUUHJpvf
O9P78k7Z7eZKb5jQQo3P5zsMDdVYHdXzMzplXmGOpzkRJxniUua7CguRZ1kGVufqTnS2eTdkNTZV
+elXDEIDVQlKDZ6rfmdGVz38Q+Wrq2+JGIvj04ttxp1FNIJhJTNT82JMVfLGMgopkJm5aTBBXaOT
93lEjHlkufpIQfSr/F07H/OSnYfS8dSy0GknE7etShGiQ4kf4c/Vyvp5qb2uU/4jv2P26dOwx7ge
6Zeg0xrAyZEUNAkx6DWW+sm03hKTpuPdVfH2kE5gY10oHg6hBdy5KJV6JfXvBvqQzFyu8Ex1nIJH
f6hlFHHmZOm+ymYnyzptp3z4lX/DUa4KESj094zN5VeK/U3BiwQ9dyTkGgir32pY/kTnEZAf89Ia
pQNMlITVetYUstLTQeZUBJ4CArJwMzHHlL/6KglJ7M+hzupwd/TT80a31BgMu9uqnuavS/WquWAp
VITyXofOyiS1RYokjNZC+XjcjuRlddVptYf3dghCUuWVXVdOgDm0GptuiCtq6ARyBydQBe9dPnkC
ylNs3DsEYkImqPJwVia0FvTP80OQru3sT1rUuo/hnfTQO0EGB4dIwgbLU8ZkJYEn51OX/7Sl7bfz
y1bfQ8MWCntE78WYdZ1Qtl7KDwTXTnHnX7E9FoC0NqrpL4R7XOZka9FADyxdQ+oGpUfboS+NLa5/
dU4fSX+VNx7jVidwSS0C6O6cztaKOC0PC8+GfeLfqL7HC14+AHHnyPuTlEwBSSj5c/X/i1WzE6bh
/QzGzyYgwSee5CzjHUeNhjFa5YrwJUN9KZaiFR7nHGlYzSFU44otPSfW3Kh/ZysiLWEHQdc6T1PZ
KeaiiWadacUpqRLk3PlwvDaEHI2yCgfdQOKYqdNMT/eUZ9DqXV2lMMQvVzKhiHw9HUu+x3TaapLP
+HL2aQfqL/SmrHZne2ExJIAhaVjVrA3tRR1VTGz7xMf3D99NoyS1P6AMAvYWzIpyaMhbG4cPQ6yW
eLHcQAr5H/jltBDHtFwMVbwcPUEfwPLFHcTkrPmM73sou0StrOVc75L2UOWcJFvCO9QFQuW5xhrp
WmKHCPQdiSNraBBGYFEnwKJ+pW1MiflCMEko97063PR7VveZsGLG6gb+QQupCbLqhrI8rRUfOsa2
+8CwKjHOGFAToH/BV2RnCWLuZP2YKiObfDiUHwdgsdj2blY7smT6XcSrHw1iMqPJtihohK/hLb9q
2CoeqKf7MPQiRCu4IWVDVzz1Z2A7oDNJHiiQ3QRQwfAdsHcHyBz+dLDWO41cuyuAAHU0fbz7a0Gc
3CfV23gDXiy15GtwWcXQbMQ7neCSsSQCC+QM6jNmyiIa1hKlgobFT4Y/8VtsGtCiY0i8zfBstvKp
yO+Ro1bwFWTvuAjX1I8XPiZnqg8OfNFnoQ8u1j38vNPzIru5/tSZtqpRXdCR8xvMLWDTbLXTwQNu
X23Eg7BOxcHAtgEWThsrkfoARuUZ3rvOOQZ6SEIPY5oiUxGsXDSYpa/X2SkGNpqOoMFov3J12JAO
9jVB5E0fweV4GbG/FX6Bbab7fRiuRZn95adrutikwKmLZovG1GNphEIXlVP+6bZZe4/74SkcKQj4
0euIMJmIvDN9gIJSC+cYnJ0DbSF8Rhnq+O4ewzK+mYUBOKz3kl+WZ0l4O3niDwQ6hxgMGP7J5WNH
hlVtPZFXJOHSv9yklOUS8ke+7yTtn9ttvPyYG6o/SDSrHmVlyhsgw70n4mi7DC9sLsk3+eGd+0ZS
e6stD+gEgRJ/lDMRxeTDWttmAvankZsEl2qr/2Z+6Bx6OXELlNtohLvRzpP/AoJmVe5QVGF/dJkU
Uwagb88VNvIxiDQqgcl95/lVWlQJv/d8+VWXHANpuN/P21ysUhIJxrk8ITeP7z52CjROlcqYF4/9
kRv9k8JdXxLrp56Ag98eYb7d2BSMMv0PNxJ9fMPa9ou5FC4tI+OjAoKa0djYN4dG39ax1LDPdYUo
9Sa77Q6Mx4Pco8EdLlWj5ZfG9rtAvrG1D6uZMXzKQg0gbdUFk5yapLETN7BFJyFhJj7XfpD2S5rz
pCd3vsNpTwSWZNuwYaI0l0AVy491vd2YldOFCpCsx5f8UhroG860U6GTwDsYWRsR9TgIVNH27yb0
d+/0OVtQ0vVFiUYoDItMH8RqEbEd3tHThV24EBfdrBbB1ZCNf8Su0DmXRsAYsrS11X1Hlkur7syc
Q99uI5uIMceBmFhn2uvPJK+F4H5JS1i6jGsqAO/AauDmCKvYO0kZ2gHAX3fYl7d5jdSDGXiNOCeO
GF89cGdvXjQiHPX23r3jVgB1i8GUTJGoaY0TFE2Tptt4e8z7kJ3yuWJkhKzjoQQW4s9t4O+tXNds
0VPEdMdSafaa++gAzHDiSPcrmf7P9IurRCfTu4PSLTZGUr47H8gP+0+QzjWS4bxZamjL++pnyKsO
nPDaPaTmJSdHkk+waLu/ziNqPwYtoe+jPn5e7mRJdWGP+Rtc+gTbDzcPAvTCZZUuYlcMLguEmqOZ
FuXdvMQ3QaWtQxtzAZ2mOeHLEDbeFjGkcAgfDpEBk53n9QTgecFt8zzh/5bXkX/PvCqBF1MdOmLW
b7Lwo0u7P8VHooWc16GN2UT6jPkvRvTF+ubvLL3peLKYBXh52gqXpzs1ybkiXS3mGQz9oXBiMqwM
E5MNDrL1lcbeIckBNV1uzqxlH3E9lZtfeBi8Gr7eA4HooPt5EW9pnmJ6mtz+SKCFrvDouGhZ0kIg
sZtrO4cHpOvwbxobpDvMAC/BYHKe2HBrB1+CCEY+8v7/ovRjLh1FnAxCP60efA6HfP4AJG7r5ney
HDi1UIEENLydgD5qn2Z+M/ZP5zyxjHDrjd5SiorT3NJw5mewq6nbHjqqcGSgnT+n2BzA2QkemcQ/
EPh2R+7Mw5mow9scLI7d+uis4BD5/HYrQzfS0vVgsSfFBh2QejJty2suy0ucUJtCl3u7PlswyYoP
kBbljIOjmIW0kKMQSwB8v6Ck83AmgJECBqKo5kh5SkrorjNsHeYr2tCCtq2C/ZgkSslNJxmJuG/b
zhSMO+Gp6DFykiKfA2r3GbiCiHIK3SZ91BO6wXo0ENmJGFLL0mx39RU1OacTS3wy7XtEGSB/HZpw
LkbvGDpV2Sdsr6k2j6+rIdG1XJNveb+xcic4Z8hMLtmM1Xd1iIGSIs7QUw1PxkxRU1yjb4gpoSuT
6Jr+Tv2A6Y7qF0Bzmzvzg7rRILRg+EjHqDqnUsh4/kdeCXh+itJNp5dYND8pqCJ/E0CIFnzboVRq
3VhbvbIi1XbJEN3IyxH1nqN+Z46dH+MG3SK3zXn5j8KaPwXBbQxpbqvg8Ed2+pbYBm5BroMQaJm+
fy3zKpWFEkpkcenN1PkVhN9/9jQpPWRy2flvwB+RCQ2XRzFfdpMJ7Aa3XURjJSEFtO8PPgSUGYHS
ywFaW7E3UhN8drHeeHwNpzV8IPNyxwIqNmOK/6jFU9PdjA6pn5zZt3GV2FJezDt6NwSK8E+dFNgX
+1nEqAi5vwN6uVOg+eeG33/PFfze7miThV7Lwl07Dnfr0ryecWilLVYsYSW+cAOSD7cW3bAj+roi
lBWGf4h3KWyaWzcpPCYw7jDIsrJgrdYUJu/9Ofwsbn0vt5CbPcFFrDpvEZlRAGhv6taT6TMZ124a
LbI1jCzMUN2f+Nz8EWfLd394O1dEVv4asP7bAijnB/QEmUdOnYeVArSsMhVEs+cR+Te9UnSLQp/1
Zkd5WEsUMuIMoGUg1OtFOzxZqgBUc9thJQXNi5k+94Q/HI18CreZOvw7OOTDJnDsmrM3+pFhPIum
bl1CR9+hXbJKxQCjIdo3I6zjqsg6rRQ+O/OHa4BoKB5z5zTT4SJ8CqCQsTlalLa3oXQ38tbgtCnH
LowYzdTmtusZbn0bwnqCkARsmpp0bQQKcn+YKITHtcQ/U96oz5Or5O2tSkcMH3WsFox6KsbaI3JV
ZFhLD2j+ImZEOPIJExyTbzrVjrIFZK6Yr0LMiHapiUDxvbO/Nr/S4AzZf2uUe9Lv0n7ut3jmDkY2
ON5+iqHyWs/xoFi/3Ca4lCKuUrSNRJQGTaoo3nNESh/YW/aaNDVe24LUBo7dVZHNPPT6p1UgezRo
An4HaA228EVChoPunjookzPNcEhRg4+wJvZq5ftRFr+OU3MV/uVVMNxFgda/RkwHZVACEv2tlXrS
owStgJXNuOm58URbRenSisrYm5l9w0JDGofNg5gRiJy86mSsJPj15M1TX2xcFiNA1BlXhpWQybr0
EjBARQ//YLogXl5B7nZeM8feMSZ0LewYAetLxRoTfJgE5OD3ZHFjbvyRGOeXTmUO7cg8gaVrGWaW
R2Zzwtu0LgTf0rqffJwRzXanelHyuLLzp2Hb5B5G3O2jzCKDUKdSRReG+wpBcybVLjtWs/F6jiOV
ZGREn6xc+MDgnW72e4ZpjfdGDqOfMlmrHZwe/CBl/QByvjRUYtNdoe6lO0MNufPUhvqYkvjZ9Ysy
9pR+McJYWQW/cI06bynHmbXBv2sAAL00pgTGPR8h3T5+Nwk7dhPVHKlkcXrNE5z2XbmdtbRkb/CG
VhbdrRZEIkNEWxPrAvZJpizAihnCqBvnM7z32ZCnkuz4Zr7+eWOEaSqghVErWAEqsef5vsLXblFR
/Yp1benxceIuIJfYude6sqDEN8AkUrQgLL4cu24U8jxXmtn0AxCZJ5C9hWH6cQT+Pwey/YAsd6hH
NeIgDmrU2b4JuW7ndlsWnvOEFyDKeA4+P7eg9TVxf92X68af68N5i2tB+jA1v8R84p1U3JMTAIAI
TMYS16GoPUCQs4QqzODTUeLNZYRyG27fSP66i0uenhBpb2bxEfDC5eo0tjk0eLqwqem2DXPlx8xs
TlWp/Xu0s9xHQAC56leJc85ltqsL85+MM+Tx/H82T8nqqWhZBa51beLQC/C7KerLelyy7LlHQL5K
YDR4e6iFrmBu8OAlmqcrO2mBU/0tyAkHTvGPIBGuoqAVeEiAGcxQD1hf8M9j27i6IGC62TIl1KKd
GxvXkbuwOsON4pKPAdiRf1o23kxCITNCFpd2rfFc0/sr0XjFJJdQNxfCQHy+e+gxRceFfHt8/veb
deAmO68joYSNXxsApHEJu42HWi/pehLKaxrhWCdWBs2JyFrnSrdq2OvsxNaFTSQDoV3XKGPrBkoc
zUs8cj3qj5Py+pt49Noyco1uQxr/9Sec3jJqWFioNwO58y1fa3ZAP55nctZ3/qhoJh3SZEw2SWRq
88gy+SMEMgGUZkFPI7O9Hny/ecxQrdhzjuVvd/QaCcGVtj7yMS5f7/Jbu3KrFylhNEb8062vCg5k
HM9hmK2yYYRuofTvrWIM9ITSaAwvpbBUCEpDwKQFuPZUnUXZ2wUVWqaMz03Z0lMEzPfA7gBA1i4s
BnQSN/T42z3MNIGE3GH8xNzFskqwK4kg6x8917+fMTJ4ID6EzmpnuqbBZWREdrlnmnnTlMckCT2s
BcazZ+AflszWIWNX2eKa2gjqTJaxKsB1L14I/r9PI47l1QhmfOpTeA3pf72RJxX8RxylZU5rbNlr
ke7PBiCM6QlUmYEOqXz2o16iPKUWFzx22h6XECIuvU8cvY2h9WTb9036QkNZMuGijUmeGk95VxA2
CnZuOzGCeh7nCRagLZhLOYoiwYslxGgJ6OXxP8Be1+XOa7iWPDu1AxWwIiuUzfHTGmxwlvmfz8Kf
EhPE+ePTbZrWX8RCeKqbLe4m49OjRwhhEut/JZvKYvU2slM35XZdupZH+25nbYjqN3LqQixiZB36
Ipdvs2MspZmkJNf86yyXJNU4++qEvisPWtcpr0775+uOeepaOz3WTRNrNDZSiFhi0pobfqTQXHXS
wdlCeDJK1ipdYkoix2tkAJH+YHh2gjCMIYWueGY7EI6bh4J3oR1FeW2Obc3dHqQVRaMUvymPhmJ+
E9nGcaHmPIM0q6pr2dwEj/Ns03kOAfnjTWKNYzEtCjH7/8GivDc//3Ida2UYL5vQFNDil6QoPOUV
oRnZVKHQr3M/n9AMXvugSG3Q+AXTrn2aZ0l0Bf9Ll4rPVXbl9PIe/0JiSYsT876OfKakuSyzSZns
ahQApHR17Y97ekpQK7estgOCgFRnZzBxo75A3SP3Wm/O1nZf4+8jfUrF4IDNRpvpb1ExjYV+xG6c
C2dyXIRavak+BLdBU68k/J6NM1jJVHKUuyeGqO0w6LtdONKsIpuU85ka5HiH2ScAamciZqGfH3bD
zekAmZk84YSExhTAHKJbLqjUeDy5a14fqws3iKmKVwKRe2qYNozZop/uNDVSkrNoZk9H12NHx2vq
BmhdYN7GUdyf7CNulcPAzZKv1Lt4G/pFMWCsEX8YfMqodQrYHPIsMYRDl6MvgUzJ5KcoEPyZXQsJ
Vby4Su+jdP3UW0W2YiKmmRIOFwV2vZdaR7y4++vk989Ekvxiuj5eSLOAYrYQoyNmkDMXer6nP5No
1X4UjURbodrUSDmfgcR2MuEsi6pBTZWruWUJljuM4ITmtXQ3a9yMhXipimdMvGk7utHKd2KqXTFB
WrVKl0CiJqVoVKZfwpzBq1lBy0H3wxnflfEJQVsavSdP4HTXNI8Fnw+WgGjn1Q4HGOx62Rwa9fbu
OMBdU/E+xRI0HRUJQlgbZGLYIGzM2pZXeXfUzRcn4yXFu0JCY/Am31JNcIFMgbypSFD/ng1HmXd7
cCS1FUJ3YmWUGN0tYmVqgzvXu+v89x1FJ3gFNV1EyXyLV76sczq8qKBkdo1kpxIDvrHVScJasTA3
c/iIVMcsRovyzCnR7ST11V3irtFo7VdFvKNaKuMb0zaLqpQt1W6tAr9UsCrySm7N3s2N0T2nMjqL
CkOrSemfTuCMihOQ9Qit2rnZ3Jclk/4lWGTu1wGSH6Q3YAm1FQRyCR1oM68aTeZnL4+HkW+Bv2Ay
54QmR1qRJJwsDmrEbXU0ZNSudhWuw4o8+NNFsMQtKntRo7zGRiAt6meBWkMNIshwMr40fruKJUdp
k4dM8eQI480RwSljsP3vB79L4uy3xRTriKKB8HVwFbOSWU4VXNKS+IDwaC6Ei2bly29d09ck51O1
VT+xGp1n+G4xHzM/jxUpV0/dHyVS4iSIdT6IBSBRoIf7CrACgtNTDOWwi9DToXg00FCeTTIZdYmv
pc12Remk6QddW0JqnfxyKctd1DbJgeUTWX0X/JhLuP4Om9QBUDaQjUoP9/FwhCnSOFXH0uCy/4jR
oNaUFrYW5C3Mvwrhcu2tl/1ThuCFwhvvZOsZvEFZ0JMBMquHLm38/jxaI2D8fFOWrZu/L3NG3a3g
VIWyaj86bHU8FZkF+1gdHACo+lAix43qk4+mVwbGp/1gH5e3IJ7oe0Jn0QE951gp2/Hjej9IMuJ2
6hAS6/ZZXzbfNEz/STm5rKa9HwhLy4ZOXzFzkp4SsUrHCknFK17y39W60OmF7FD4PRMnTSMN2IBK
POtYplj3pzae4LYVqS8goKM+p5fhA/4dpmLg2YxU/bp5d3ZKQ9D83E66InmLO1bMAse0EgHJ9jhz
Pyk+Oa32x4WA2vib8rJYmUgvdp+HNK0+jCvSTql6x9AC9kEASSXPcK2zqaSNOlnKquP2mO24wyub
vpXdm/aAqpOOwPyquAYehf/UMEJt50dl394l/3fL5tgre+rCtkgdIaHCwIpypTc4+U3w280IhG4R
9tBQzGduSU1EAR4xKjmgwicbERtF3UP8UG3TaGLLUeHjlAD81sBs5davd087gqsdScTbBcHk38rn
SxZsbIpG4HKU4/tnIIgQpOit0jl3zU/NmkH+wdOBYSbmZe0ps42zLaGnnLRYYsTIYG9cQHevElI9
mUpvkZYhwtYjuR/bQgOr6aWFWSYDtODs+hvd4kU/NauYY921xwKrvbSTuvd+j9EREVlEGhwTO5z2
F5dNrYdrH9dTpua8mVXwt9/w9nwnZM2XSaI0nMJ3ikTnAlHZFZ6LvXBrqL7g3DwM4PVIRvHwV9sM
V3pJojX49Wffl9OLmTowYoBLbIxqMQlMMeLhzzx1eYMcTa8Bpj3d+R0xwkNmpj4p1sTbYNMgvYpD
tTzZ0XqY9N2Y7N5GUtPjU0MG7RVv5wQs1+Qk7Kbyu/EdywTCIANM0NzWoneqUThEYOVWXwRMpbuu
cy7z+VD3cYDIoM/jowXiHQz9AljBJmkywmj5Klj1Och5y16ZPFKIpy6NP87w1Yi42hQ3IEZuf8Ki
Lxb9YiydnON2xgo2dGdJxmWOpP1TLg7qIx92KEh6wGK1Hi0pJDoFLRBmOFin7UFJwZeSaKL7MOzS
ruwTtvcL/ykYqh2vlBLA4CYR4JHWv7K9co5P8EK+lNpxvShxQJ4iNPWsVWBUHVxZEuR4s6xlrA7g
0b5ak+mCwTRDrCntUYzoqNHSsavbk1O3+yaZhmKB3nXCO1BzTNnjsU0RPJqTYGG2kQmJKjD44CPb
c5c1R9Desm45qsET76U0aPdUUOOmnny5tpdVROWCe2E6qgXwx+XghjvV7GFFzl/qws5wzS08w3Ji
t/5LMsEQ4k7BrlUdYWK++dJl0+cV2+pmlOMTFj5PkH3NJMiB1o/rq+kJbV9QP4WmIcLwAh0BFJv9
niv14AU0yf+8Xj21uCp3MHnsQXrB7qQLNfQQefDQIKHVDEx+HUshTpgD1AyRUbAgTZBhk0R0XkK2
CpaRoQ0+6AKfX8PNVw9vCy1u5nBTNdrqMOOu7wMSkdYtiFk1BLk3mGWCsWXC7wVeiam2DluI/LTm
S9jC1yzQtKZwpsMKGNuWir8RQJYf8hnaqiHCOg5gcTa8gz9HCm6zSjGC0qlUPCa0tPpl9f9TDTRd
SRrBqIiIsCUrqgkt+H9yFA74QgXsKIJTaLHAm5Lmkn52vVr5ekHPCU4mpHSCMTPR8oE1ljXgP/74
ebf2TAViispid9yOO5EOL0Q0qWE8eNxUyl4C+LTpOWTPmsWLoAHHG4Dc+DmuVtAGXBB3rZA2Uj7P
Rji+uN0vdOMng91PW+kc37su9XV3OvKMDzWimQ1qW9b8mMtOq8ffn7V4m4QlYRVqPItXOopGvjOR
gUbNddCObszcuQMjD4QfZ7CHcUIOkk4eAhG6PfZHXPzZk9TlzVH8K2D1n6BE8sOqz7ew4Gl/tSxe
qZSNu8BtR4NjMlMhWu0OMH5vOxZJS7HrFBZzStUIEzXBdSMPeKn7RgDY9a+MzjWiVKzm1eT7Bq09
QpteUMmPSC12nU8qKyZE0gCpvvGJmjex/MC2unpes9M3OuYQ/9qv8rwbC2C413WQt6wpJhcJgqXp
UYM9/gE29lQ7IVRI5Xk4idFenyosRtEuMx9xGeiSASz1qAKLq9yvvdQ4NjwNlJ+iyGzDYbao86mT
DVWeHysWhMk59gWOH+yqLw1ChoanP0BLXQojNCzUiePHQSBqAG+wIXm56jhMzmtkEF6pt1SuZdXy
7JcLAtSyojkTJ5PM1DaGBq5ES+5llQ+ngqDfoecU7VfcFhFycv+3zLsegGyQ5qpWczCXBXma17l4
gkiuj4eBJssNWJbxaIae05hUrPXGe+Syc3XECoXMHvUHSn8UFj1qCWadIA3NDjnf/1B2/JERv5S5
/FrFyFAGt57yVAVIwIfq30bifv/cMHLQE9gKdsqqWwl2QA36hkCgYxlLeaK9Vg1NB03WtkV+J/7t
SKxoX04OolC/Z4m09aPBVFapHyDYfX+08EPhalohJep2CL0t81YmNnxHLRAilYM1eKRavFJ7bsbW
MohuSNU7j4KqqK82nv5i8Bx5WLcKFCzJX12LeVu3rLZLHYTY/XnDnjJbclC493L87vj19LBS6tWn
sdEAiBo/3fDnUkPcNiBTT3RF4Viae9qnbI4nKXm5CxAOwyhwoN9DXL2Zjrlr5QIjDCfcFEXFw3Sl
dAdQyaT5vSmb/J0ARGslURs3fGWwyADjsh/4oiq+zS5pVWZy7MkY3NDsFdgSKf068Vt/LTBpIBWs
aVghzUn59OwYe210hfcyOE0a9QRZoV9cn53VUbnojOd0gAGScY3IHUyMJJ90XWuZgiOdChrBaXix
sCB6BlMAKu9/w3D0m4XsNxt7JqXKVXiZIQcRuLvqhu/SAXivh0q3SuJbePoTwDFY3rN9VFSDbbVV
BdXZan3/m/jfq5jkiN0ibM+FDHKuWvZhYZN446Q5NIuH6UJj7MS3/oNwsPB4sMtgXbPOnezZITgT
e6TXPwFN3CFOQwp8irFLXTcm/8AtdQQ1bNjuW78xQlwSqojHZDvKwOaU1eWBKNCtEGjLaDbnXYSe
JOxKrTToSRCFf1TwcvSvRPeqitJ9I02mrWBdZyngcgfs/gitg2LrpnzlhxVs7js2KWWOlmizlv8F
zRIHEKUZgqtjesUHGazc9u24FeiqUWGQeyQMcAy5DBAvhYrEKv1d1t4c/U2D6/1lIQpFjvmVWJxw
Idks/V0DUXZIUdnyZ045b+MF0uycTGeePRoHpRA79SitjGgYPgs8dRwIuI/BQij+P3JI1S9F8PNt
bcQXRNoPN17q9KbWIzrvodl1lKru1XjAGCn5hGuxywqcJS7RZi52anB5lJ9AQ2bRD/Eml7T+qLaw
I96CiavfeB0xrD6wx53hrrxyxYETJLuqstq5ifal5pDeNptvVo2dLh9GH00CjCiQOT4w7JnSzVrj
/VQ5NX1qNYdsbjaazWX9RNGW6PfrEa6xsG5t7CACvEgkj4XHexOGoMlHmkXWFAJE8mJ2Cnz0Xx2Q
jL4pNyBSugp1aSj3P3EuynyEUdWZAij5iwOARvtkTAcFxEAtnYLdYh5d2tTvuNgCUjGjp607FTMa
LGsEnmtbTaqEF5OfTqxMb85S2cX9+3f/R/8kGP+nc54INcuaYNiAGPpPGrQIocEsyrjV7mi94FEG
XEeRu0wgsN7gstsbjP/zFP3G43ATYabsYR53iu4RJGoT7gTttfqcT3cq4lZ3ZnAgnhZYGixLfSnS
ensc2jrM+TuzL+QX5GXNVUVHXh55ZHGpx3XOx/0I9pc6xB8jwYTcPJ08ogDLKg1H3UbIe5vYSNfl
ACasDAfE/3EdgOGWNBQNy0mfHFptB2qvMfCK1sc+yMmpfoXvF12xPTBhg2d2dYqHFC8GNbE6XjBg
CkhQhBLtnvh8PiJniAXYFnu2+RZ+b7gfiI9ZRF5JJEHelijNu/UxykkRnn5fnkyrlwmpwpNpEAL+
wDlRmL6x2DcPRwDC5Q0ALBXx4tADFScADxHS5av2fcTSL4vxotRsFzZfEUlP1otdA8FJmERyJka3
G8X0ZRARBS6H8TCANYVxQ8x/DAjOB/VDgdhpPaC3ZuszUHwdA6NAguJk9cfxAGPKiH1pHb3Lz5cl
kRXIqkgrJD65r5L0IAhGQdpd52wVsFn8ytAoNFZU4OGkE8jZtdhFwS4Fi0CNmogtHL4EGgzTedj+
x+/VEbSer89rRyZCRALtJpj2xbofWPLWus0lSQgRbWB79XhgyPWxJJtmy7S8Lk+yD3fyF7Uor18w
aB28VTfCU3vYMQLQpichRLRvHG4XMEwcjvtJyGOY2pgry4r7QiNjdlOr4W9VsaIsNVRSwGuSXB63
S/cyVonkbH5EwXvlwhcWFMJFHq0mZIoHTfPjOQW/6ghuNT8uG777OWWDdMMm7YhIalIPr1OV3qds
1R9yDcbBd0MyMoJ2tjCHWjUC88yCrOpFPc2E0tMTDjUJmgeoZfgAWZ6jkAkLzdmleV9239VasrOI
tCqe5Tgx93Jd9tpcJz48ipyqx85ZUIaWWSa4pqa2TP6IRVtQYrkj4j572DMVGQclO2oXPwENoC1N
3ts8lcFX5Aa/tFYrNxJsJ0ksCUFEbF3/zzk7WJ0zg6zNj9pxVH15t7WIRj6W9zrl9r3dPDDGxLbR
zY5K5I3vI+0p3DMW5aKwwTJvvYR0EmDcwjxgNVu87a8lGDYse//LwKNVEjPKHvZiDte6+V4O0UhM
t07Rk6NjK+LfBWLzvONsMoHrCeDD+DnTZ0jPU1n7d4M+Ecg8Mp+LABRr168/D+TZH+KAWGvtE1Ml
SfJMDDH1ZzFDKqWhdJ2DStwXygwkCwB7jEKrfjc//9/+E8W7+F+9bLelJO+TVCeRhV/MMIWIaIxj
M+HAq0cXae8SEmoe0OiIjFVR0tftWKBZOEm0/7xP+wcTso3BN4rf9rgJTYaYMPzWcBgV3w3VS2pw
6+f/ku8VFGCSRGuwWnJErYjzqwubRluzjW3Mo09lB6fQWf0/aKPQaCPkjjYDAhkZLbyK++uz5P0Q
zj3QWuIYGiKeudavONVtAPlIgZKueYA6xN+4LFCOu2x0er9FF/p5dnI4+Ai+TlOMlDMZPnDGVnTZ
tDOt17GqZv4RPKjF5R2UnljnY7XQvKWbhiMcLgON2y8P2XWB3nEi6wYiISC2Yxgm88HTJ3eL9pCw
Kh4EFhn6Tk6WEk2ngskIWmHl+/N96WaKEQWJ+/GZoKxzWX/73gbLaNJoFV96hms64J+jDb2yu7zU
Xbu7YW2OP23BDkr6aB8DSLIgXdd6W9KpX5NrDNoLt1u1cF/AJOiednceFCJP9SpILsfmwsHZYJuV
bTuh5btFe8rxfOrevtnb9T5fiWPkuDA6PzovLmW5322dhdL7p8QqyWNaQ5QhEujt6af+QR4rAChk
Y7Yb1RHyr56VqieM3SZ+dwADz72h9HSQ647/LV+fp+fe2ni1+K8oTOOAl79w7Tj08yGsZqtDUJCi
PVYqJTNjpYxkYctxqDVg4++ARFxJl2IDmM8GNsxtFAUsFsDsTOOyiNoccnvRSBHq5Upt3IkTal/S
j9ATNdhuFStRDjHw9unF2YmirVHDpOwGfaEtBbr1jDnoyYos3ccRrfbWcfDOADomNDX5U/FwoXvE
ZThxBEDqaLmG6nONPqNhfBE1yuGEDsJ+Zv0XgWR/qswZbtqzQWoRepiK6jGpleJ+KgGrklyYKS4m
6Zeft7OPyPBfHQbPMcG8uPPauUVJeHZBoBliyj5MaPKrKGKfaXOed23rhLh5Sd2JsohwFlNOvM7X
jO3eYmWLWykg9ityaupFJaD9iAoaL/+0keYYf4JiLWmNNodHm8NaLsp5TfQW3FgyOczkoBi1j+eX
t+OtsK56WFn0CWCK4rC4RUe2nCG4+4s9dy07mS+DEMYdUWLwTdu4Uqn4ux7B2Hf9JZezIUNttegC
Ebx9OazCF2YdKRT0Fwm2gIw/OcKEv18mabmaOPf38Yq/QWo1BFRo2da/CLHArxoVmgkuccczxAaN
gqiqLWnu/kwZs8NDRaAye3Syn4Y3U4frBj+n25iX0ZQ0Ai/oUG2b6aQbuijCOFB7JF11Duh8SxJ9
i7Z4c+IGDgCoiI37CN60OJoF6Pj/01mhYKxiCCJ25Ka4vaSly7xv5sdPIJ1qynNDUIBFsitu6m0/
era7DXz8KCUhPaApsq84TdY8RqxpG0W7Z2vOWRZ9PttzWfPN9lCwMRygWUWyAaMPIpkxNxfPJqYW
mOM/2J21jP9VZG4PaQLpuH3TAI/JomcRm9IH1kPo1U9dRo4pVb9oGAC13unKbtzlK7SxEfTpF/3r
lss8D/hyXgZV+tSj0aZ96Hi5UDhfC+R1Z6nmzp0AfcMUMccQ/FhtuD2sXJqhtDLM7SYAniZGEI6o
B0Fk2YJVXCZJ5+zYbfHElY5p2qXyq0Cplh2IhL3t8P9HLUWdA7FvVlMnMpF+JOkiDgSid8WIpflC
3Lo67Z28C9Sqh+uIMEFeoWMu3jRHxV+kUAYvIpIqAe3506cqIb0Mpi1mSjlEYnZ93QHQDZSLOqk9
/TjM354UwBj+gTvS98BMEpKXi1h7QfM9EW09dmDjSX+CHIaAg8ZXLGFcQ2nVS0YYnmiFxZjWlpri
ZMf5iDQuxTXHTTSWyI9oWXh2o/BzprVLCVSMJxducbXMiJuMq+ipDtOxbjhavF0mFPXLNApsmhr1
4zvk/SohDxnKNgTMiE/lZSYYFF/YFYp/wz0A0v6yXRIHped0OgTvK2Ks1I3yDNXbBYJ/XwwuYmpt
M+/CKg0ELYnBp8PKUvdYDhZi86ZpY5+VSa0F/S349G3pf7Bgi4UbLCb56FM8vMeWyLR7beckeKUM
UUpzy/snltiJtS4XqCw+kq4SPG93ixjdQmnGYvtBuj3JcIYrB6nAuocfBQ2tVuT29+dTPY2WwDKt
hGcpGjlcNoEZFT7H/M9JrbG5ic4O0d+cSpApoQUKpdGbbwLqMFL5x5DKZ1I7nb2jn3b5Wtuo+u/H
ZUfrct3N/O8pL5jzpTU+5i61z/27alxCoI4L9ZcPa0W6MLLlV4ibLhLy4LG3c78UP1gWWYIce2E0
dgy7zp/wW49DG01tlUlS0b+xiKXLkTs4UggPoVFsd0yOEdi6B+rTxOwBGVVuzWafEZaO5ZxE/YHO
w0rkaog+NOOmQsjmS+qhHIYvSNHwy/lWdbwou1Zv/pE2ewqx0o2U507QTdADiFUTngMPn9/qmUyQ
a4csL8Vv4nirI/VybavhQg8HA9f22khJHWYUrlswH/P4zYIy9QRXhoaDMTqmejGVAwER0coa8s6T
sd4tv/jH+sPONQITZeGSa3cjMhN8z5TxhLKsmCJcmyaluG88kEJKyV7BfZfCVn9JFBuoy1Jb9ZqV
uYwHpKUniAmAsG4gBoV4PSkbk+Bl5pscMbYzqbNt0LgHd3W9QPQ+Cgo5stutBL6arwa97ghYRNPn
zSq9hAzKlDYBNfuUjdFG1z6gxPeskqlg+hdToYKNTLWCrnAGxgVCuVJFPKJANZlDWhennU5xbcAy
elwzJVYr3vyPP8d5DDcD31+Ttj1cfjFQLdzOT5Wmq3uiwDyWVzc32zeQoUtE29QsJthYXD8w812G
HZ0QmheCd8Rr0Z9i5rlzycFTjrdXEFP1uifJd1bnnXumhfJw1+f/2VF43dp2sOK+qVTK46e16oBX
ObMLF7AdqBJzCztvb+97bss1IHVcAAmy8nAok5KBkzzZNTAOtPVCrFWvq7atIwgOFJApecFCud94
47on+BHehN7/9CBGl9+YjelqT1G6uBf7sBJlS4S0UyXov/kUkMufkdsOUrUIGr6GbyW7EMKSH5sj
mtBhBvHTrlmpbt6TfIrwmcQXLVx1XsMFQPLozMtojta+FwiOEAgK8/bVGs2P7IPpo9OZh9wHKDmQ
dM3G1mLryxxSMbvJQwkUYFMYaSkkftxWDVu7Qa/ITNIhHDunKiHSYgu6zWvV35Noe5iL59otVJgZ
sNyVMCP7zrPCSkroKSSHBPQG4Z3kJ2BnXJT7jsUgx1TVBOEDUhOssoU9ANAjdxNTthWcYsVq8atb
nKTM9AmMqGfT72AjGmTBaCzXbK2keTAaNmFtCoC2GA4tIv8oWF+vmDNMzSkQlpBKDoL7uigBHDqN
w9IeOrdvetnc/gDW2U7u8n86y4uDvkvHnwSOBiGikBv3GC5ylq84AAnh/DGdjqDgUlaiEjXQrBYc
1IyCqC1+kPBAaC2nJ2PqRaiP3xV7ojy31KHobRmSu7Huw+zjP30gCCVx1KH8yomU9qmD5jA0kctY
hkFzGHUXX0DkjcSd9hJcK2nzm2Ja4IZ3eWnXqg30VxDTxNs5F9NZs+IJmllFafNmRWXwAn/vHnZt
HjrFLaU3WjPadQ0Re/P1S7/TNDG+XFoGZi+I2Xd6PKTBQfiOQc1quhp05Nuxg//LNBfxhc2g9EM8
hmesl4HnSNHfngnEvHuUfOA42zyM8JdPpdibr0dE/VNfsdVclVmkBdvkz0N3cVERSWQZRurX4SLX
R3vNlE1CHeYZuiUFifSJqAWJRZ1J+GFYJDRHBBfwnuzJutYPEzlWk2LBcphmnDLx1IVWo6mR2lK/
AM4SFDm94C8YKJihACCNdtJEVzSpiNP38bR/FBv7tUgxbT0/OP75WYgsjFMUyMcdSlxSSNnhhWFa
beFUn/O1KL4AIgBxrMKWrilluJHmDCW4W5O/fosKRLYe+oy/+pMEJeu77VcoJKo/26AmKJniEmpi
Cc7Kdq9TpLNh64/6w0jxvaXvIHJMTax3hWCKWAGtLLBMCJ24X1gJfdMHnI8jfr1M/Xdl4fLWkd0y
S1GFEaPw6GySfBWt9qqrojcqJ4i6cvxodElRyBAEoead8YI6v2pfAi9vOQZD99OopOgX7ynPpsrw
d8nc2MXdBt4e4h3KNbNAAMuBdi11C/QPyAzql1CnL6vgs64mV5fz9WXQigRbrnRQ5E901PqmpmY8
iLmwhNAIKqjdcWP87t5MkBd8gqgf5pSTd9e93sCZOn+rvthfZKnhETVY3PnGlGuSmJdEq2Nu0893
k1ggZwKOkGtChXKfU89wd2fv/KT/nXhITtGxViTQms/SrLo9kD8zhTlEv91sK+nzJGt3ETLY3U2n
UNEWT8zaia8kLg2WE+lJaCpUnhlJKOMIg6jXVAUxFSCItD5UJGK+vSrjJ6+IWt0Tqp+HJrMlSA4B
Mgy3xxrvsG9a4fuY/Rfz+77QTGzP+XZcemSjyvdxKsZGEMabDt2RDi9o/2XAezRaqbWSRmGJ/hgX
tZFD4JkNR/+Fe3ivIuV/tuYsYrBtNSv1t0b47jIETwnYZ11AKId+/HoXfjOZZ8mYv997iBfup2iE
0zpNg/9y7eyrSib9AG+qHm7TkdiHaiu0nKhOQUosFhut6UPOqk8sVH6FFIs0JlLln8kNDOC20kWs
kZWvxy+un0ac+sU1xNKfv6zmQwHi6WVCA8Am8uIP2H7BsaCDQ7U0VDwhIq7E2RHGpUULhZfuwqFG
3IXXbouc3IM6wI8XcHKNnQMQhKfAuk2MRUCnrGZnwdMJdsvQHVckvyT4ShV9IzA41o0uOSlCy/dK
SAEW8yaAJfpVOZWxhfac5ZugcPez8rP8HHpQXarPxeoe1nxh30W761s5TCZbBvykw1XOdHdg3Jul
P2V+yX3cFThd0s8BdJFB65K98j3j3uND4F+uLKina9ZvoTsP7Jizh4LtupkN2jM0+LF8IimyPSUC
bwN81YcluMHvldZGJwvF+AMH2J/euWjseyDacztTGyFz4GrfnhcMovSjcC5zsbbUb+RKb1Dm0Lll
FQFNhq08ee/A9VVb/yMTM8IcMfE+pbiKkg2VSRTNCcbPF3PFKdY2VSf2dt0rojR98kv79NZ10i56
UBaIM698bcRn8tKtgp+saL6t0tTCD0JHoh+8bEVEXx4XqP5Tn3S18JvMzgqRM3nOPlXWQnkZjiJF
46lmPd/4VawPerWRKL8PPDxMqD5oz50JfXTknZsG9E2rVNS+xyND2tc1IE+R9BANnjMPumj+l2MB
Vey9OpkwlgSrYJCaTM8ev+FfW3vcl4EfU9smSOKMdWhhB0vpiMBG3SDBZK1M6N3/Z7G/d479bJJd
QOk4XDt3nADCAT27bbdcUTZ0+IC7vKNGyJENUiynvklxsKsr4xJ0tgvHfvBAOLkSw3E6w1gAkvwi
/N0wxWbH3s5PWo9lvOGTtPyoJH/NSWGWU12+GIzzYsW6fdF+0rkHht0T4acbYF93tYUufCCCqt4E
wGDvZW24Wfoe1uf75PYr3x+U7f+dReAxg3SZiw3TwkhznUj3uv8fzbRUoWwRVt0WQByQ3cIOCyff
m1nEHENrHiYtVtsz5i+HK999vVmfYBEQTuJSUp26x3ROiw+wUj/AfDXJ5Ox+L1rSIvOnfsYmb8Gi
xOAxYOyaBVIHwxRLKbPXvSgU0pn4j1Z4cgbfwjGxxFCcKx7ByvyDgkrwCkrceAnsmRKEnvULwPuP
4pjw+p+w3LmWePJMRO53N6Hq1hCX81aBa9twj6VwJPZxksGCLVP1x5otvkx7mFuaxS24/yLcNuJ1
itUCmPjSW/lUPt542UwymVB5oSfECP2mkFCLn22uZZQ+2YnCE74S6P8RyHvUrG2tv/fVwMXJfZ+c
wm5i5Lzo4GRfkw2B4ZcO+LCwAGx927b3MKx6GdxhkXpX7n5GBJYuhiP05ileGe+eOxysPwNp0OSr
MtVaLtBAy3dRg36zHgWMzjLHKSsCiajhTtlwP+CWA971PuqdWVqwN81b//+eVoyikMIWE8nv13Lx
m+rJOcEYeLXIY9rLkufVH4jesxzTW+3NM1tyi7uRfaSD/aDoaiXCAXznh1V4+y5pAV7UH8UmFEey
BjfNVfUhT/a5X0fwdcB4625M4sCic4dr2OWhckqNj6n1FoTzGwt9fT4cHADr0oqPdz/ZcotrULaP
57PbwlDQxNU2HrNpY78MQDNtchGchrSy9ImMlbjdlyR6PCgIGVPHnwvmQYqdJCG4D0dqCX9CQmCJ
jkZfgisUzSo/ZYixj7s1vPwiJIvnKA8nWx8rSDpK0kNT3yLvGaCPHpeS5x+f3Hq7YVYwEalk9fXF
pmsYE50FfkhpDe5ZiFytITRTuQuikFEd8J94FA0+Q639joD+426A3GRz5qXk12dyrjn5A/B5KzhX
QSYSo2kCdbES2I1I8zHAehpuIbM24nD115mUJv6jF7uBcTCizvEWowuSENSUoK0cP/ZyEdHLhuUa
aDJWmmgC4o8Tqnzoznw49OFZkxZBRyuv6Jmg/SwBA1obqmPJ+Rc469dGXDEKiAdLcMqFoZT7UAxy
MTrNiZNdI5ZDww5/PdmETxaZQLw7d8FxjJikDp5FlmRqHzcfuOOpezvkOMgCKVPUdx3u9SKayFVA
v04cfI6BPBD2mbcFr0sZI5xGPw0q2WjBj0Z9RPFlHurAvfosVRiy/98t2Jbj6w7Io5egul9/RbdS
OKYWhow11aUCmfUnA5owNL1/NhKQ8CeZV5D19UOOqQLCSWpRpdTFM2YSANTrkdrArCIaz5q1cezV
mS7Bomg78Ys/QjS93CVpUHHJJKZQis8JHSGIBie9pxgDtaxlQCBRanTU6RfEqIUUxO8JTYNTfBDR
DItNvDwFAAe0IiRTh9OV+x4la5IaWOtxUK7TEThUkSPRPZz618F37oPV7HbpSdFhqygC54jITmSu
d9ZQ3fdRnn+BeCrEtkMvwnwhLtwMve0/8zkyK3iZU8umxuGOb5Mvew0f4fT9tYKYHyJEPkOPMVYS
n2avK6xC3/+Kp0mnFO+cbkfLWVS6GhGP3LMgJSDG7SUlBvBSv4829VWFOr1AfoVFvMpb09g4wZ2X
uRgqO0eTIua+FwFr0n4IDeqi0BpF8pa/DbrIhur36ZUD/a4I8NWWT+3thtFF6GWqKZTqSL0Upp0r
PLqFdiDTyPMvsWhpVGBfxh9/QS9b8jnnheuCzcjJgoopXUqvgXPV7irN2ND/4silxP3Odg/hjsXL
1Ifd+PAo0w0ncLhYrh9Yb28onwCitNO17FNRFg2+rJIjcslbdIgfNs+1LJKb+k37ExUQzme/qSzn
i+hjV/VasYqYcnlzQs9kJIVbxyrk18RwwVan/k09w7zOkMC5/rGWSgQ4y6vu97LtXvxa9cW9sfNM
Bl6myYJatJzqbR6W6fH3j7UCgMRUNKILWglTFT15pKq3ADE08s1+S3MG0zoQ1yHE32wj0gKPcY+q
wFLgxVFK4njR9cX1LAQC7b0+ypOuYQ2JoOVG7agPdQEZrHjKzW4bFwoVt2TvBYo12nZv7A5OhEVG
yNHCWuGmBEYbJ29ksM/nsv6J+GO32sXqidKM3tIoRdOp/T3Q/sS1piD2H7VGFNnI1uQvzuKwK8ri
nera2JJRIpmOfg+MNE7n5fY9mrbFuYYstExhRJIrB7U96iFuXlmBLyPmJUXY/iLXRKCjLDM38BW0
J+bFTDvK0PGWwI5IRLYQ5MlXmddFzUOlLRXHvM4+9sTjkWOqVPltT/RjYY/vk5qjivO9fYMr/kim
BclRTydNyW7ax+s28jv/J3nSycMxR2j/MNzVzNf5RrBsNZooQriHd5ry/qgOuUnEaLt69QCca6U5
rWP3Gdvum+k46Ac0IQyQkqmHdd/zke23jNBu/xnN3yIs//cyV1mCvHYxr7pSJrp85bD7MdRdSukU
EToh7E2PfNycxlCh75DzJXdYtAVHqPvCQgkNQK+iznwJEnOpk+3t/Zgt+WxghLxlOpCXNngvVY18
x4Zjpe5JHJtjoJaY2i4YHj5dXkCV6m06BWtpwvC/FUH+Uns8gdstJs6kdtG4tsxC1jhjZRoicVnW
KqMmjbdr07PaPLu3mHRBBDWL8X6e/GSn2qJkaPb/jrOAalCRoodMhwnTD70v6sfGmaqgsYLfJMj2
ah04uU8QRrFSgArMcctnQnVvwKeBWhEZrW+ovNOw1ywvtQeeV0amGtUcVWv1Zt93Exh3kXgdd4IA
/xxzWYBmgNfbJ9SB0YRTHGD6rnRZMeR5zu3bDApSSJLJK8U55Wqx8AeKTr/nxS6osqvdSRkUOG7f
WF5ARMtTFt1us4DEnhU0QbIvtP8qqO1det/YnNEsXjsajsu9y4ESgMWyY0vJz3Or/Oa0PLR0iO/s
nnoGjpKEztcg30f2zTd6bD4WuqmJ3eUhPEHB3A5I1QtTTZ2bELa0F4JjXk7F/Eskp7WhFl4FOnPC
HiR/hZsCILNOW3NRHJP5IjYSfqv5XPwiWwgQXp/NHl62eysxjt+HgPjQxv6tDg7ICj8SNT+qemfA
HfQsTv9SHNHDaGwH5enTBEGLoN8qkSev9tutY0KwWdTRnCimIwGi8INrkAotXumrd5Xs31Z7K6qJ
5F2zvII+ZSJWfBzzdiUVRNooiQcWSCPbDaJrfUKzu5LyXMmKlpNHeIoa1gqs/gacVly7cLRmhLMZ
t9VFu8vGl1nSDtSrK0uO1ElB7BoYx4x4vu0yenfoJ4i5RzlWqiX6GkFJaxKp1I9EnNquadK9l6B4
NYvcIYq4m01nneyMycAg2Frf07ccur1IXQfJY5LPIMBjqOo3gy03SgV3uIbN0DowMvs5xdB87828
5AVbgInyKM36mADgqW337ablnLgeKDxQvkCanQ==
`protect end_protected

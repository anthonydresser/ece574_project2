`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fqR67s8cBy/jbTeN196DpIBrWP6p4S7KSN05JgotCa3DCQok9PHpESJ+/YLHnMMyfVgYu3wMYulS
KP/HOuKOPw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o2f3dkiR8+1URrsaFkNAXM8HKCsrRh7Sklc6YYRJzdPn803OFcwNwVYhAiEMEOIJg1X2/T1BTFui
EQHVCIO1VCJStauI6Q8S2fTEfSbCGGuhlpfWUvhI0fluVmKgzRXGSxAPfzqyEe5IOj2rwzAzUH+w
I3b+vGSxoVxUbGLho4o=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ad3ngiL9tir1+ET0s4S3c+66wahwIoOVYNaNS7rfCSvbfk2aPsU2XB63og9D1Bg2SAX2HS1BQP3j
tM8/wIjLaDyunyJe0pY3Vy/MM/fpwDOYJVu9969hFmFD+MKjWmgclI/zBXndfn3HroxBNJ5YqbWw
T15thS0zDy/kMUmQm5Hhk2FofTiKZfDwJV8qMOs+IPoHxa32u/A5H/GAlLbYSj3iKXMDwdX1qvMx
Y/wH/Wca8f1dMVlyNgkzE7heSVl+umU4imcINE9Qacy9ksyf46mM/SkHQVg8M9UEek35LLEeFt+I
FDFYvl4xwj9zXwa6o3hy3BjN/8PdN/dXT3nHmg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
17s30izSWEvAAgQv6Vh1FDrqsfTI6ntDPxRKHcyQC5iftYo778GlTYz8H+ZoqnbRpo4Rx9iJh9p+
faDV0wcwXzKoFudL9jIBKm+gYqfFEvkVVJxOAlF/jWjG2nF/VmEXgcx03HwRaHCNUzX7tGZCK7Sm
cgQAO//GQtSMc3uUvyg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ru/nQZrQMQoFSUTnxErYixiyU4ARIhOaWewtUIoITFUVgG9z+gMss2pnsjU/kUZ9RWEI12+FXVka
+gRYtVpCxIPUEsXDftLv17WDI1tjcj5fWaceTamezhm6KUczosnGz9+NwbFG5z/2igcDAy6nQkqh
V58et0XyT53zqrn13mIfMOozEcd9PQwsZNuQCbg9wSERwoxnPdBLEg5UXNHZ0s6ahlbNehvtbbgl
yyf6RAnPelMgF4kT2YNl8xE5TPA5Ftff9vYHl3maAuj8YQ9wGLdONKEnZno1f+5yR5ljo2CbWnO+
oSovhdK1JX9QEbIkJ2QqxqDve6XKaLZUt7uHvQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NF2iKYemPHtuWn5hnoRCuPNs4c5eCM1mW9ddVILQydQ1OxFb70v0HA+tFCvBdEc/Oo23RE7HCPKv
BmrL9RcO1vKsdu91oZA6FdC/0KF7Iok4N8JN7IggHYwqedBTXbT1G79t+dcJQCYpp8IWyrFodnmv
7En+ptUiWn4gmkvJxLwkJl9miXUxtGBSTbY+MIpFl4u1hjtD6y8qRkjkITWWniMoIGON3+ShxVdH
vJ4+gC14V0VTb16Wd+kS1JZLUjkak6YQE2Y/wI+gM1SfXQv61yNCkzn4q8Fc5HhMXu8wvrAjPOoS
ZjZwz52Ph+N3YHEMsKW1FO0on8vy3THenmVVnQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 59568)
`protect data_block
pa/mXep56TnCuXj5k+7cDZsyudF/BgySsJRGxM0CTQyXaSNE43YiJ69HEvLxTJm8Ea4pTJ1v9WXi
nTRcVg9K3DHOhOIzICKejreObn6KOMYE3ly/M7H+fhzllYOKD5pkvsu4Ux1JnnXHSlhOWSUZUS7c
akygS3sF56u1cIP9LsmT3kOOiB8C20Ky79k0MLRzdKyMX5CNfDaZY/+5/DlZbEinHEAYlgI+ubhf
1+JHzUoW/aYf+ivlEXVCGzhUDTLOi1SemQRP3R6eadXrxH4wowmWng3XG+rt5B6A+2pEVhkvXiuv
nwQQBrpoaeVML4tQluMXwQymGOluh6vygPPJzCV3mNcyJk8r8V2ma7/E0l1iVIQ+/QstvOlEI4dq
bhgc4ypBpyqv4HZl4wZt3HzkpHk+LHTuaSI5RFInUCGElavX49VeGg66jCNfi4h0eKoEaJ+snOUv
Cdfpn+jy8/fR0sqSvdykRXo24Oi04CsiiFsTO21vqKIETnWoUzil9E3mRSe4HGLTRL4/Q3d/Xxd9
dPecU4PJoF/qKSx225w3yONkXpONYFTkjXh2SQOGY7kY/xJB+354v8/faGuBw08+01XQjvlfeu8L
Jr2hWT2QnLOIwBq5fIBc6FbGf/HjseCm1m9wG+fBDvSUL30NOPPrhI4qYWLaiZMkjN6QNkppTcZV
HEyxkuc2zEugyBQBCWN1CLTHAr3RTPyEeG9jAe4NQ4tzsLi98LfBhLqT0AC1Bb0ED8s3tgUgrcyo
+dpXfFpHr4FkcbD+as09mmyzhcYiGj+H/fujL9Obu8uz/NVnc8yXKidI6vEN2JQyVQSJHIhejbqe
Bwz+YblQFaFb3VVEoyHOI5ED/+XEspIMEBkSDpYCnDB11DUvMK3VITT2xE15fSrjUMuURvMrkILg
97tJ6ZreA8Z9KzBIu5A4VVXBduI6mIHslV09aLK8mELsByMN2Qq9XMBPaRiH6KmCQ+UKf80VMdxx
TGz6iSyvFhRRhBsEj40ch1X8EjY4MqS4gvv5+K+Zew5IbDw0aCHymAC2AmR4QneS3hCzFPu7PBPN
e7GIPnyi1LgrDCGvdvemFQN6btu0krlbV4y74r6cyP2BMkDF9RCItZolRMIFmaxDotMWa4Vp0KFI
KLZjczrCwXW8qQc62hAnB233bkmA2MMmpUxWxYZy6Nl+3wn1FrCaaDIK/fOKLdHqX3boWNoYwlUo
aQ1BmDNa8VVAGn3HrtgWOGHeAC4Y2o+WBLAUqzI19FQw333xAE7PkAJmg347xHqVWHkDYA1H/QZX
twWAb2DeGgvh4/GuRFuOCKWG+JTU4pHa9pLirBParpRlpr4rswbROkhiD/G+suKBDgHODtYxnbOI
LceHSRYrA0amKpsAT+oVSepr6SOGc5PWz719S5A0o/IYwU20i7U1zcBYqLLJHh6bOJZj5hyVvn+6
D69YK0E++fBcKtUlKXyNYPeIFujHn4RGbP++IniBGSPeujNp69A25jEdu5v3a68v6dBnKGw85O24
GE+Rzf8sh7MsLcjDR4i5ju+Mkgh2UiRJ89MVdM7KqsMs2sXwnWiFx24z2Lb09jvGE2DDGlJEXZqH
Gd3SiZZiUqM7zM+TrNse8peYS608joObRsQfkJGi/MCMUogc6NEavUUTJySL2HgeKt+XE7r3eq42
p4105c9Xe2ctgwMNRH4y4Ye63A+vztyMkooQZ3dZkQEx8vPlU3WJbEpKHYD6eEP0r+0Y1vaHfQFi
gykPngDmfP6VPuIm854uiDhmpm803PchsU6fOIvv0siq2xfNLmS332Fksc/EhbrYlOjQHiIVM07c
ryppgs5O3N0MJkepzpcQ+QN8wBSV4WbcfvKOncI+Lfiurn8zIEEA7wo7V6Wfbr6M/FEyBNu/iJxB
3mcLY/rYLBqWxXnYAuzygj4UIxvd7w88Rx0xj4ikwIAL10+4EB7iHJb0D7g+Wz89LvSYBeGhwRoI
KfEL+f1RD8FREqI2IUC19tP8Wp1aUWWcRcpBErrFd4nO4fRFdyAHs24Q9xLpBnJglL9Pm7A8aLpO
0bCehNwN0TNMLNrCt/x9zN2ni6HjflH0IT4X/Hv/F9y4qYFc2lkPT2Qmu9Y811KemKDtd3ZGYb81
DA5ycm1vFUiL8MmAx6shSOP+TQd+bvMIMCbj0V+y55jGBOS+zWJEDuZ/vRMRsQBx/35sHAEyCzyA
JAHVbrqznahmSPXHiDGCBHn9+SX+8WK4Y4JBPdZBcBl4vow4U8F7ByTSX5xXh8oRbYwqrcvCQAjT
wlZYnPqr1UuKISqgrV64C+przm2POv6BXUS5ggP4GU5PPrhuQ2Al29abMaVQL14NusizApKWl29z
MuHDRTIRSg3Xq+IGP3rouURHT78zsdGGRTY6HAgWQT7wZ4zpV1zg0onlN0dKPhKrNUQ7+snKjdus
r2VEzXA9Fr63D3tVU53rwKl6Ds9Ksh14+WqlwQxmSYgJPLXVJbHvYkLLfL096LjezhGvMN5QDkAY
Cd5Sd+OLG+TaIH06bPMx4eRRllPaY8q6/IAf/n76cP3g52Wj7eZAUFuNWc1ih5GTC4OccG7UCCDL
UvwRg/ijyuPeE5GxnlxzEN+WQUsaHqiV4Zrkpk093Nq0uEyrXDI0oKatyff75/4NJXjwqHLZ9RLd
BswxK9ntofx8FYJM1Z8mipmcqoVfZ1f5y9V8xOFPQn7D5nA97E90XRBHQG0LeUPtESFmWZy4kZzf
IvNR9NQM8QN47FTLwiEsXl6zcGwknoTPxuoTzQMCLrIcu7kiAZbCGynaKJB1M3fWQeFG2kHTzGX9
4CEG11iWptElTnRibzlTQStEBTXqPmKQgVXhsPJzh8FrYDN4NmyFQ/s0OIj8bDkegt+DnNFMsZ+C
kICi7FEHKEtNZy+hvZmzV7bi15mgWUL+G7X1veUtujcQE+mb9cPLb4aEWIfzX+DWe6r0173kkLUy
aCgt4uzGyPcwdS/fEB9pBKO3cl5aBCbz7DQfGHZfj+U0ghjP6YpPtFg4LltI68ZBWrXdBV5EoW5H
mS1yDwcpI+mR46B8+U1BvXFj4cv/2DZ+jaya8H2kvnxffX7qFgYElKd0rS9RDrwrB//pa8eV4ucl
Y5b8OFj41ee+r1O+DpZDX/ziBfFG3fR5Qvjyfg1SBF4RxEdfNZ5dRKKkKrj9ENuo0ij/rl58+0++
XIV2NT83T0ahtxHd6M0C89mz/MgUGZugcI8aRKpNW0uBxS+oMAyEJCYAVnva4SAQmnLuq7qU+Q4D
+7y/371GyI7hIp/+xPMnI6VlLlnMmFAb1AcbdAib5f4Pd6gJar7vtVBa0GOKTgYC+fjAJz3uLz83
nnmXo1Us1TKJYx6mWXoqd3GsliylNWE4uOL3IzlvUWx/LMKgjrQhD5bB/nE+VR6c3uWdppoInwJU
97VoLV4JLeTFOh7dJmpUq8xHkTE+SwuLtUTz9HgvEIHQ8k5qN+RaNAx7yCNSXx+B1/QhLZ+pJ2Ws
9XLgSPEoMFa5TliFLMCkYhBHT9AZ/eLhtxYZiaFXNhz0JR2kIsjCa7ldd4I4AvD/ZWJy+uNh+50V
6fZ/ktFgdVIwE/9sPgGOKAUCU8+Iiy3NVPZMZS6kcrZtCH8c9mzscWXNnU108mJONBLNe0XRKLys
ZwDafj8SQoAEf5HaxU+8m9PmTuqS4yZgdwgvlFEuCYGzxvZbXeHTc4rxmw0WUIakDouYhipo2okN
HQb+tcGHG844sqdmuAi3Dm7kClEWAltuKP1JQlieQkTWxO2Ttdk8H9Ux7w0VACMWhAzDmsqVvuA9
mcC45ANehZEHK4X1UuRnGMcszU0BUBYC9jmQ5LAv6EmyYN2KjhAoCocW10IQWaySTdfSFo7BreO9
tFHJmVt214yxC3L2XGcYGM66MRM8oXP6sbrK9PJ9gGVw83pPxG8uUdXi5ocDePH5kjyztiuFOPcc
4OiHbP7L5k371AequshCgbLrVQwV/qUTU8qyiAnGVSyPRuPtLz4nid3ogDwhVQ3XDyYy1VctfoOK
tBRWqvGiiHG9qC+peHtpwwyrF0MQ6RROGCbvasDQhdmYlodfOe79b7zCN8RxriiNl1bbhW0RCntC
T/jVmeGIIYpocd2aZyvAUjVYRDQWl29LXfDBTB5ixsVG/dGO3ItfnypT6xEm625acoBnSZiUtm4q
B3pF+K1M45cZYa6C3bpXXS+gJcKu2mRRzhG+FjgAX0CVKas0oUZoDAR1i8Qap8lH/ahevRrVqeuq
JD7QCc0ieUFdlQjcE2a9lH9PhfcApyeaBgh9yNqDiJzNBD2/Yr8So+BGEgdBhveujt+oJrkrBeXE
eQwxyXS8rLSWKMsaQDO706CITsr2LRfaQTT7i7eAYZwL33rxABbeBfQgbVVlKwBF+IlMWQ62feUt
m1obRorq05/4xT8pfR/iuCK05E3z66ULuzQvoFCoGG3Y8RrPFjGPnaSFDGmQRYWfrULIDDrJsDj3
z6CE0sXKnj+K70f10Km9qEGILOftFd8inl7oGweY7MeuGwkK/Vk08xPf2lDa2ZY5XmXLDqqSPABM
AJNTcMRDgJs5MMSZRRACJyyZgW2LsRd35JdP87h8vbA0VRzBzXpmNJIxLjd3hKsYKlRq2uxyuwNv
f5QqA1Y/iqdfB0haLqU2V+ZivYhQCtL4kqPx7lztjtxGLFpwS/m6ch7g9nyZMJoYCJTFygVuX2im
D39RESODGEKV+ru5CdWjaAMEJSwoZXRxjXMRqq+cCtLaosnns8zgUFOAn9n07n8P1xuNeykGMz+1
150oc7tUvDJhDeB+6huo8ZuBiRyKDHtS4EcCHf/yJiNm/de7ET0tYHPqUo3+cRxt/srm01QK3RFe
9eBJ7/zTRUIiXfBUAxIGQYr+wap43SLCf0zI+exJrRW9DxezExUt43/RxP58KS9u0tyRtaMytqqe
KevONWJwnd3PjOZhp6KME/v+ATTPVj0/a/eTbBLNx9yeAvqtsxxMT+whnW5doDEea0xJutPA/QKK
OPykyRLlfQyX0iUQWvvw1GUCLYkgslFi5lG31D+lx3125/PvzElOpgUPT0IuHpQy2qWCRUg+Xn78
D6iLBXo8UU/noisdSPyx4C7yQwZa44S309inVd2gVBferRGQu4OHn9+rC5nt1rWbz+cSID+rg7Jx
6xdXlxpnm3mU6NoFSaG00F+ihi3UqSfPvzCQecK0C91yuD8KwAUpd1aFTG95OWxDkmySn4k7O4Ut
k+5FlYKKBLrvpgKd3vTec+DUvh9zl2Ce7qR0Uq+qxR/69IC2IKZo/OnITCeMEFRxzGUscBWaa2Cz
nGhYOZu4Dq8RF8+zwftfHBYW427cf4F22gBcaDXq9T+i4psQFIaZ45NyjSnYdeazYafTTWcPQLDL
IFx7zPtO0sw1M+cHAO7ZvSch5/MC84ERgtwzVHRGEqYJIfe46ok4JvUfZ7e4z8OIvsBYUltyjQFo
3zxcl0Q/7DYnmEq3fxF8BXsPAuBOMAKxBU6L54AqJizBPRcvEriZe7aWs6wk0NhiIaokGQ68bMaU
iKJNf9iBI6ds/RSg2qLjgxe0UZB6I1KPq6hb2XROhnDX4njwkqEJc9u3qCYheVExywpdj4BYshHP
KwubQT79xnOwu0tN9TuNGs9ZDfRvVY4Nlcs8QqA8k1RPsFb0fxjzy07BHCLw4jXYwS+jQ0/KgWJ/
ghq4PuWE8QKH9TTcfJjiOJMUMcIhDZLW46WLAI6IkxY3ciKm+skZE00v+auR7RvaEYr051JYB7Dh
wmGwnyPum/sEaEVQPs5LB4E+dDDyOPHaegyfWCoZ85G+NV3KDIt3DhT9juJVaVN0zf4iw6q223bq
VoCssi38thE+Ri18bIT2TIpNsl3+83kp/MHwn8IAh98L9Y93jWTfLPD3cjLQYRT3lyiPCht6p45F
KGiAOisro0GugSiBHUAUVzAmBS5Ve43EtJWiMGO6rGu4blDlOmvzh1tPtuxreup0NvmL85SAgyP9
1MdTbrTetAFjNCHSe43e8eg454Ki/4vFIecjgUCeIOC/1OtMZhktK/HYVgFwzJBSmcF8Q78SguCB
gZINt2xjqsEfuhxZG2u/ZXbojVe/S7VfBT/3k4waTq7B3nO7OvvKUjOjR94iWp4b9nWq75t/HtFM
RzJHYBVQRjq9LLrSKW50VHsq1wq6OIger0xZ5kIGihdZzPa3T+ETcbyBOYN2PjqV+PeSFxd+enAI
viB8vJu3iKtMDsV9QUth2MyoMBbteZPixbK4QksKkAd3mdb9xZRP8Da90dwe4m6a/I6FhQ0ndzIC
LzsAoT+M/L4btkuIAup0eWlgvK2FJEYxa+18103f9IzKxUdDlALLTLDgdXefVqXxAaPJfYsHPJ2u
YQuRzXxzI3fkuhaqJ4zRvAeLGpAbgreRVhmQYyS+iiPnY2G101FD+ptejqkQVnrsOZwWPOrDpTDy
y5t6SzgSbk4asbXYktVfd7/v2B73jWckoGKQJ+N6OdP5UO8V736p24+FgaA8Ac79G3qww8bf8la7
KyOLW6YPVDIxxchikXDLoffDO3lydODdNL7PF8D4DTmQKTLgCjFGLK3699Chspef6BB34mjnMavV
7BPpv+3iqN96BgT6S3c2IrEQ6Xhlf38SAvisUds6os5ogXg22uwD9jjc8RavRMZbe3iQ7mWr70zA
fVflk3ulvGI+8ewiMoMJgUWOHOm63HHqC2w1Iq8QATFMUGos7ZVSPIiE7r9CIc1obN8wmXEZvKJ3
nMBmtwegbj/vEA+M9LhElLcRfywzjcerwh3P6Y65hSqjF5nR9IYE1Gx0RnR1gO2Vm7lEiej1I5KQ
uJUKwYCC8Vzdpjz7JREIb8MkhLKkwGDAJ+2Xf0ljigcJFsamFBWO32cR9QF2VXHe0U/rS9V/BKR1
0dz8+tYnuG7OKXQQg/HzBA3L0DiIx/8cmYt2gUWLrSWXzWICoLN5rPoPkOqdLuTbcrdynxkbB+km
WngjJDoFbEuH7ENPLZ9yhf/3ptXLdWbib6SM5RTxuLv6SLH6lbxjA8DG8ZSCH/kD3HF4e4/+fq1X
iCdvW1RqnIUJ5VqiYD0wilUg+AVklSJ3y2zjmNAiqO3osm4HdTdHvtiCdpkFzNYfT0WjpkRE5GoD
vbmBKMtIOyWjbxaa81AjJvmKdEvTYAh9on/1Y2D3QlQOg1fU+WJKu6Zxuh6+1xzGDyEewqGAACKO
wAdVF9Hhb0UQFp2AneAl5tPBSE6QBIVZ+jXvHUgZa36PgoJk0mJmofOMX4zoBxR0sHJM+u/1GXce
3FXsn/AgMtlNT+7dAajOQaA2NG3R3cJAZ8QFlBWeLVbAjDNw9P9Ec8HiWi7zigTvmBlhDM/LbxZr
4gBg37nde3WAikNXlICGCPu0wfGXUhdNSiyp21BQfMiflN2DBAcbnxEaZhfT0zN6/0zjETmIJ5jA
IdxOuotGq2vZ0dPH1b248MZBkxy5X7txdQYi75909ur4besYWsXsgmLPuu1lAko/ZfZDrJ7IvTN0
ete+OhsYjW76d+FJWQncEmNH6q3Dg8XCoQMesp7mf+bRVXfJ7NyNJQWZ3DhLk1p5xqfSS0F2NrND
uDgONtVpCkyQxWtKsIV/igJpV1OIO3zNIpfM4ahHt3PCj3AVsaKTG+KyrtQ60qdMrWQ3Ps17NmlI
uPsMzhSMK18L0goN6Er5tEhB/I6hA00JrrhXKYOrH0D8uQuXm2ntNfotoeHeDAsBuykxn4+FBNGe
xBfIbqbg/tM/m8f3kc2eWzjALkMc9srowUOGzUGQAfyy2xlV4W/634NavKZp2XjjmWnMxbz+06ZR
0X5b4tnoTYGBqLzn1+eoTmAnLcqivXHYoqC85ye1g3qyf9CTVY5uFD2OPHwcejt/tHkKpIiVJ1+3
uBtjgDFHnlEDbj2e1FINck8OwIWU1Kq1dpsQcq6pv1SRguJz9y0J8b7af8YL9uFpKpdxNDtUi3zc
viI+2aEQfHwWqrWjbY9okrfjGbt6Vq1zfgblaeAqmvgktSU9T0pIMi+4hNWjMYkrpwvrtXmZeAug
0bx6okyS5X2hjPTAZUghYQhN0tUVG9NWx9LQAbnmjEiiCOENL+5bZKxwU8T9r3zrXxoPrrGT56x2
bW+PdojQ3u7CJSdTeurT2CcNMyvzs8xj/vN+TWbrVQyT0zXsXjXI9lSnPf7LJjdLEoGV4fP1Y8RD
j19Vg7e7wn9CtzpdRG68alYgX4MXdj3s8+NvRB5IqP5nv0QnKuJ9Dkr+bfyOohj8R1VHo4QWexQ3
Z0YUoNoPa+FoqpJuQ6ZbqbjA27o5Qq28w+gz5rAs6G/NSe25Ac1dJv6pIEi0rpegQjyrB5nKky65
5MzueRwafDojBALFRC4ff64Z5Lev0f97sHaJfHDXVoU5umGrKexrd2oqz8bF9BwEHk1fPW6tvoXb
gmvpO7xiy6t4699pDNqScDTh/43Xeb4dlLOrKKAvweymJaGV9S9iIBx4dOyreknGNI7Dk83bv35i
VZd3fBhg19538Dnfa8QOzFK8xzbcc014LZdBjoiiHE540tXsNvho4asCio6eK9Sqxw8qj+5Ezcbc
500/txs2cYS6R3DqcMP2BrVC3/xb7WWWH76vKNGqRjoQVpKV+mnq+vzTE4o3b/GGp7yPfDHDiyjn
qEFhxXnFNHw7CHPdEzZMfVXu4AFl9KDL8xfhUjKU5iZkZaJxKhPYYzkzWlEqEfPrg9iv09DWwLZr
048Ji78uCU0ErqRGfotg92hLL2ggULfzyL6v8h5g5PofZu+LZNkLu+HaKIeDGDedYZpfLY6EInGr
ic8XoC69oFMRK/nJLthGA+8amDmCGM2cy2RoTSY57zX0m2Q4hQTfk1BHgswyk3/WsWCqUYq4ZNIP
ygmUfwB7mpO9/8Bk5MByBz7TZz2gT7KOtaD82Zrs7RVSEy8T3cVkgQZ41gEjLNbeK52UeI8Nqbku
HQW4HOAXK9/ysfPbDO6DQc+wJsxuxAN8tZfqbbNlL0rsdDsvMk49f4oRJH9wg8Qwo8L1mi3YY4EI
XQTV9acZHqBzaLH+6Plb4PpY+jLZUjw3jI6uh/48XnYSqh/DIaDG6U6XCiSviF4XQgrfJCt45wty
FpSx/iVMKKk0d3OwkMZDxZvz8OgE7BmbOS6VzIl8excmIATYDgvRYohvSMXJuAD4zbUj+afLC/sd
yvJlcOtBjEMO/ujZG1RcxNomu4TuDYuuRJROp2+sS/0gAu5uJg0IJ6wE1f1YJ6WyF6nad2r1w0St
RHqbVQIXQgIqEpNlrtCmvguAHv3iXoyuHADIetY0rDBAPYiwnqIcstRyPFbHbhyyE1KzdOnu0NqW
IPfo3hLc0xIfckC4pllzZ+j9fLnD6O88SqELqf3fPUu11VHLtMZICT6qTPA6W20pmV6tkNDu0Dh5
2nFPcADAsBlzQi9eBqJN3q+A8L/kexiUCekrM8MZy2BZZAE+8M1TD4igdhkSJA9BoM824fujrzEX
zkFkus4BYF2/GmzTWJQy4UTSTMCKX+1b6L3OneQabvnzWD9j/1+eXyfOBhWVgmcVn7I4zQPX6laX
XA5U4xbAMIFOPEcG4pTzH4U/OWEXzxJzfsEgJ9vopWz4+Kv3CBzhvGyXBaN+Q0fleBWbLe1I8VmT
GJGaDUgAB1NtqnHdl/BbgkHhXHgf8v9yXeHEUFg54Hh2JFic6tlb2Vc8lU87avpppuXoM1oWzM/T
YPi6zlwtxhNqUQLXLKoetIMkaX55ou7hMGtlXSeIFelqYrU5WGfg30YQsUU8fEAEDI+PWrd/5FdE
vXLdoTJ8v4EHi+Z/XmRUh8yVqoGY+daGX34FU+Sirij2y40TkQK2HF2VbDl1vm3g9CYcc4AGjf5C
8tT998zpeXYF7gvdp7Dick4itabvmOUZP24v52KMRINkTi1l4/CU2eR+nk9jPnpm0yONJ6Mr0yhO
tMkwGf0ATZ7AJMm0wV736CJyyr6fGtjG/KyG7t8bXg2GjyzXvVqir1Rbkt4t8flHvs03MUR9DpGv
XKbpaEfLWdjMYwrvlow3YmMWAqGjLhAbOC4/wpJY0aQWvxtK8sZ8A5jNa0OpHpr+WpXGSkKGrEQ3
j+cAwH+9DJag17zcLDAPWzlcYrpvkBwpatY/qR68Pn9dNOcW90RNjNsAGelbY8nusfUEdLEhfYoP
s5hckr0ig7FSh419ItuDAK5NplxEpdO3VbPxuCdcHcN5NqWnL36YiVYh1JrT1MPwqdfOm3uAVZMa
gwcuyHizs12rmg0BUQEWY2n9HtvFzCYFzzLmgXunicQlaPEBqSsnXpIGZykPSL0xP+HPirzjRtIk
Wh8wBloJAxbHq8DRT4y7W3pvo2d9CVxh1qU2yQTcpVTJnI7jWfuJO8Q+UQnCS2K5wPJNbIOa6qvj
VsnkuLlQCNRkezgYe39jnNPfhLp9sCU0+f3/w6/zZFc6Y4hMYw5krECdRVnqU6dsF31wLieGPCEK
IpXgLW4wwebt6lQu8fCDnBty3e1bvM2pu1axx00RREeRmz0qv5qZvLOzkX3HWYj8XZhOI6Z5B61t
dYiO9l9u859Fr1FZZOlDvqzXqf/i+D7pAOenvOCTnuq+GPRhxa36hRnui+Wv7RMvOoqLnf5CEAda
KRyCp/fQhI4lV8sEI3pTbHx09nd/bwwUozlEjHiKAHHIoc6T4X9pvz9o1CSRPBs+xEOxKuRe4eqB
VWO8zVEfUaUL8Pcgp7ZfNLIBa4lmneD7tk/5uNUxx3TFvTKn/vuEMpzp+cmXmhps2/FVpMq2eUJI
mZ/YxsbtBOuhCTDfv0v6XHgGa4XSd6ExhqUUEIEIkq9I4B18mDCz3q28uosu/BqJBLoEYulY7L1L
5hHevXWcaLd5knlEoAqgkDL2PWwXxcCMktSKxYwj9ZrdQkLZhBqfh78F1ZD7LFTDSzddLmugZlb0
+IL7nPqBfi+7eT3XtXz9rBEoExHR6Wez+IqqkUzD3j2hqlyeWWCzjX8/mX2Jz+tvsseRP8ocq0BB
HQBbLh8E5LntcQe5b4O505QtcdBkqn413k7zAw/Y6t6zIHynUaBEVZujdFC68lS5DcGvQCpDKufg
+ppOlZ/3SJbg243wZDPVs8oODPlDh9nJarGABiUfh7YR+waiFipU2JhtjGx/DN2WOBSvSkdI9k9Y
y+7Nkh7qEtli9+WFPz60rEALRDS2yJ41O6l2vZGXeT0tmQOhFw/DbsXLZXpui1XPWuSayywUwDXI
692b1JPFdOszf4yKb9wjVrnfqcbyhGLO/Hfpj3v4eA2M2qHLSbMQcXvljJyusFFSGI28DzbOHl9z
OXssqcZmRsAHlea2xu9AFbW+GKZw44an4Fym9jbf1mjHaKgSKREeS5NUM7QVpytx3Lth2C1Km+V9
6UNOpRzXiZ+i38qynhYZfe8bQI68IohW8YgVddEnc4t82ecK7RjON4V94ihxNUoczY7rPUn8PrHn
Bs2MeHpGwajX9MpyyGXyZvWmtKBaukPgnMTiOJnE020D+Kch8lj1q8FNqkLHLRplCrmSnj4uPMgZ
t1UXswakEqRCg6h6Yhv2vVqdRc03OgfHN21zOYsyvlr90YE+Wy1VDZZUGeBtGEh7feisuCcHcEXb
4xbZTEoLWmg8xxyc7GkjjEjIl/Dkr+iQTmMJn2yELDnsbABtiEZvOYTuWvHuHG5rbRd3mgbL4bIy
4s74+H1Kf62xN9kkF2uQ538/74/XqlWGN+Tv3uDpy1yh9I4hFID/rdpcI5E+W0UsvpLWOox7YfS/
pVD+iTVImPTXZjLS5XkcBF4FRL86Ny+OU479jHnMt7/qvHqVITW+jvoFdOdKVTsTIueTGWopmmG7
6oS7Yu9FOebTUATLa4m8wvWBK2+VTAMOkNlNNIyihSSr0/WJPmy54Ur3O1a3SfnEfMykeEmQ1M5b
TccX4AhQt1oadkcnKJDzrHgkamBJHmnof5KFZQunTuA1ftNtXib1RcAt52SaMWGgK8t7JHrf3O5Z
c779Qvry0gDx7geeouttN0nXMP3v0T8Pwz3D4nQ+5t/2sS9B5lyHX4BhIjg/TVKtrZcuIJfHRZoc
/EqaKfqzq+m7md5tofIwyKFA2dng6FqJmJYSuRzRedldU38Gx5McxaYN/P7vtqY618CRA3tTgBGo
2TL2n2BIpAGUlRV1V+cx8sk9Eum+JRHTmb2aB7HPbwhrn2jXkyBR1WaMbiUa7p3GuKrUIb7rR8rt
IEgBJ8XmF2gDUHQIl+2y7xNrnQLNrrJ53QtuNEnglO7SnJIRdpJoiYVeB3X/0mg/cAniWkOzhC0/
s4aJE5+RblrSw7bNK6gZpz0t7xQ7K6y3GpApowlZd5dnkATu1ocuEVsL/1o6CTDU8nOkw2cANJNm
39uHAmbSTo9WtMCgIWtKNKimA8pm/L1DzTzht6kOwQ9sIL5pvr9bNyUGbQDbvBDTM8qP1g9Oz1wE
gzUihtdVIgBf8PcLWWiwaM+dRKjPfkyV+8xshgqhDoEn2Z71rNkbKa6Qs0xd2/LwvCwf2CwnywyC
WXCJ1pBMj4HF8uNJEEPRnlMZ1+Zx2TEletqoT6c867Q6d38Mv/njQbwX4zh25sL/tFaaKH5nfTYQ
atkhYldmw/RWaqDwtJENfe2SI4K6Xq5TYTM9dc/L43lAxYuMLyK5JQMVj+3k+auRsdl3e9AgJjf0
t229i4AMIww33+h9ZzL8qlokf1JkjydCQtHOv/YMTSZnp7BbeRXvqRpnCwknx2p7qC6+EM+4k75F
U+l7ExD5xXyyqfPujyecheFgdS+UgGMQMlPkL5EcTkwIGhTxZ73ybFIv3mkpb9rGzvwjRVZpUhZs
aIiBnYjdSwjEcTiNoVG3IEN87pChELD643EO8NRTVxXCNNzgm47UD88/OfroJipqM7YgF/utbWEp
DCzxdKVLGnK55AaGWlmoppUuctMxi1leDFGO5t2EF9nBb5h1IqETKeidbBHVwYT3J6uTUGDP69Pi
1rP7j1EcKYaX0EiQ2dqS7G3pqNnDy8Gz88Lth1/NgNHp3MNvqOrQ8lNAv+RvEqeLGmO32hKvP5UH
eBW+hI7+xKK4U7ZSc3M3myfPY3sQ/W+/6Fi0eN2nfNIv4LSU6uzpQNH/xpSLjPWAVvZ63rozTkyo
IApIkywubQzkQN8xMRF2hx/mMyRQko89zWJxMzf4jFoFTdJfuV2bcujKyDhOlSQOmAQgUIpvDhAr
0gsDcxWvXqeeJAGiX6gyfJx3pW4pwOgimfSWbgzDoXaoBTYMHCsg+5szTdBulrks/EAkD/hO4YNz
sW8MNEbx8NRDKvnHsBNPhxo1fLG1s9Zppv6TbEAZqIO5e9IWegIgxTUTFKvYBkgXorPazk504vp+
vtGksAAkXus1gBZLOI0O/a5kbvv35SSirG0f7o77hMuxrtP6kciq/Wd6PBI09fHSKbV+7ICjK7eq
THjkwSbQKdU3kgaK5lx91aoB9EniB9Ds0EC5SxN06VUHi3ntioWNNM0bY1DVCsYbj1KJYAZCBPOv
w03RXqFds7xMirFhA7C9GZSAUoc3kgGXGQXTDwLNDqG0/r9VnlPdOg2Uwx5zJNwu2n4aPW+g36a7
R/dMC+ND4m9gtMNDo3BuoK0l2C+0rquC1v9d1ChMlJE8v9pgu5L5d2r96DnbsIlNRW3sjE9lSD2t
19sHYHfRuuIJU5w/+hMkWbJrin1oWF/XM559mAoKMsakT/NTYecsvokm4ogzE9eLkAKeZ6Rmcb+Z
6LV+iPKFPcFDsU797J6puqbeJlSrt3A5Frvig/vYbC1sXyvjH2hroZcZbeBkeiERhSEuieeAVaFz
Q1aC7iPjXO1hWBvPrJCfT9RAn8aBrHTykx77oRDm0cWMbT/vffpTiRIK7KiaWMJZvnIZVkZcjRNA
fIo1i8NPTb3PEDFog8tAteY+5JgtwobZZeLeseNBch0VK/46kr6vifbEVkWTdcApejuAhqJSMCJB
csG7EzdhbldGJBXYKV8EkG4YSxtbyiPOllfOlz2bvyt6Wp71811/3/9D+Tvyfc/0S067UTGOEKqc
EtYb1Feh0JR10XBPLzdJ0jdDyijujUNN1iVbWbKA3zES+xedPGkELXViTIdWyPuK1nD7ILGmbdp/
M61KN8DBcoqWhPz4LAo8aeh2FD511SAya+9VbUVsPb+j981lLmI3QRID1LaQ+EEIH2pl2M5u22mZ
FrjWFvATWiU9eKqm/GjQG/UtUpJqgoSnztsaIlFP0tSHxeVnhlQ7U6lJJ52r/992raeULU7Sbf3+
cTKJiLCjmr7iI3jItosvWnMet206XhqqOWhQ5GVKbwgYfQp/Di5ss7+R7H12Y79pjt5B0yp/EZfq
JfSW1lEqWGa+zkwc4UQ7D60fujVcQcWteMdRCMG1jiKO7A1+gZ75qRyI7goE4vqOpQe3ZHEe7Rm8
rP1iuNXhdTSblvEj3TOIm5pv9TGHPVGNrqjkKH4r3WHhQDHr9ITiunScEApyTQ5es+FGl3Rlf6uM
cHbcpmtQrhRkgXY0uJsCdWiRio9yk3ct1WE5Sm9ZX914g9RNA6HNQ1rjgKQPx0nq/EFH6MfLW50O
s9iL21NmuKlI7GBuxxgKAgq2QTCu/1sEJDpePSFa9jnnrW5CFkJRakomZfPWuFcYU1CWTWmwstTI
90wTCvQqNNi7/edntqfHbtypexLxntz36lTZLIaqaZT60HKmc5H1uHLuNeCAv7aZIttr0wVknLEu
X9irGBbsU8uwDzMe33+GDxBdipZrKa7K6RkCcpVwWCN/d7vcv7eplMNM4vvOCmX5/dW1Oi8B9S+X
v9dn6C+70XXCsM0+q8H6SMR48GxCbbcESj0bnoxQfGxRkSnxMYTIk0bAOEkV4Rv+mWc7Q8I4JhyH
RIsjxaJpJ93bcHGdruGj/2/kMs6TNHf/YjNB7YpXggiUz+02HHWB4rc+r97ApcxI4L3ab3L8qqpT
1y4fiX4tbOsinMCHwoiAhEkJKS6nlY3HecMc8l/vvcCV20HNl+LPjlAZ2EJct7DjW3fD9qf4n9OK
p6sa4DxHpFKido1IG9nwxMRfOYZzc0F7K2gADaj0/fE8U+KEXQQU/h0+IGcN+914I24vUIh2E2rV
mHgCUem+1DX36wspjBPi5ftcES7ZmeVL5CxNzhIZQd+vItM9yKMDf3dOXE77YQkBK+2MX1CrQvZI
BVNznHCjMRf+Pq3peaZEFD+tHAI+CLsS2vK/Pb1pH2q+7V3SQQ9FQMVMyY4PeCA5YWTEjqZ/ofq2
CGjYLNiqHRoqh9exaq1WFLS0OG4rZq3gSt6l70BXssTvqWzYljeyBsWn2DJGfuGGtm1Mo9ohn66u
qcIyJBJ7cQFPpJBhFwtAYzHPWSijXp1cBmNpiPDTXNup7ZnszJQJBOfjXLYZW3d9o8PUywcPK0ca
PES4mNtxFFol9PtR54JmwAJ2nVQALwnsZ2qYdn7Elgx9D/ZmMDaeAbIp4h/PMcBxe9i86qh4VFgf
p/9MGezSb/TU6SB/d/a0hSSZnO1hOAt2NEOg3v0k4XWa2OQBRxXNtx1JbGAA3PWpNftSvrDH54XN
L8k21y40Qc4XwgFS1RXHlhEqkcAwRsQI6WQOVQX0f6/+RyHb5jkzGrhsrAzQP+OUVosawVILdKAn
DkTn31OZLwqC07TKJXefR7Zj5lGzrQjXeAFOXEJ6yAF18U2n6DmBGvBGRX1VdUN1kRVuqVgkjCPy
CFYeZdAOwBB/m9A3WEIFl5RI41+ysTLmgnQSGTmCbzTiZ0zMgB1Pp5x7HUufBQQXoVPGZqc2pmio
zFTLr7QWL4supCgNswNv26+8KkVIw3eWCK9obifZVK5YsxaxxTVzGa8ZnfiXc7oBl7qCRaxEqJEl
ulp/bWyqWNa9a7mBHNQuE2PgVSN1NS1A9fDsDvjxnTYMC8NbAeoQMsaEjLe3UJaIY9XmmyCVA55U
vV9KEW7rT/X3WUoyZ9mSNIVVa68iIHK8kdMf9bh+kCFB5lw9wu9dkCc8kPJYY5NV3ae3XzDTiPtd
q6gTbka1H/Mb6XcajbTeeHsfZ8F9MZ7nghI74PHPw+DuwvkELGMWiu/oESNNwLwKR+mX2xrTDKc7
iEOYnTa0+56B7rrFRIgGBdplzRmVWS88n6rQM1bC5zHFk8+x9Kk5BdiJQ3UQsG70/Il+uGJXZFX/
jTynViqEbrjmyQ+Oci4n/tmnz01ZISj5hgHYs3bLV23neaARiRMztCL2n0ZC7upCsem3nsN1pvQd
DmVAjUoum5zRCFkodiMxTZdVUGwibJs7ZcmIfiSb7cskoWQdY+IxogSeCjKZp4kMm8IYljFFyelw
LDoqAYaW+onBMutr8imdQF7CW+zKOc2K9QsLx4NZLXQqo3mFgwMcpENruXzShapoe2trufgkoWqy
2/2TDoiKDJMv5Y9yg1hjAnFMKDiZFifG3yk0XUsl41t2ZID9FgMJfRF1IkkY55g5/CjXbXdg5ka2
/rsVtHbYJqH/xM95/mWoI+0s3n0+b02ruvM/0PR8LoHs+jLLykgx1pgqFLxcRue/F9rK5yp/0wq+
ULfVnYCTwrmODvmJJk5YZXTCFCvDgWC0T9UQnhPs8KrbFVmYe18VtoSRlaCzrEeIrh7A44yXo7s8
Sv8pNZ2wnskAITJZLbsqp9+2WhNgWxd7SGzvVLjwwUUzpZLcrfBj1UVRkkek7gC5Fs9msQVbe5J2
IrP57yRfKcLOisBlejdqEAsaWX2f7bcXyH6rEgHfYyiKoq7RpSU0nwjpwj/AzFygkc7IAaeHFY11
dv29/fHBtOMdWAY7S2cZ4gbhG9LO+2updkNsHZ/h69MmXQcdLNNX2l8Q1qtJimpOXF7VUo1lnsMe
qqOd3fJln5ac6BB8dEFgDpAZ8OARHanrC2UiPd4Ayqgx3QlhXn06l73dstPveqnG3/arOcq0faEy
NPNTGA2H0NnwdyQAidHI5FHC0Aty4MHadOXEHo7yI9JqaShrR9hQGnvKkt9Qw4h3yeE6XMhk3KrT
gpJD4Lg5AS6WtsTj4O3qQi2t9Yzpvzx4ucyUvqJAAeffggANsL6BqirOiYjmt5J10vip5IjK4pCc
dwCT11VwVYSymoPDY7F6QI5xT4hxRNPcWimaDHJUqkgGE+XZ2ZF4MyruSOEaWUnd0oFqUkncWv92
SbCwWwYZ714+vmgF6ev4aCu2d1qS4rjMxF+F+XaHS8NGsoOhZFLrSrDON4n3GNybwQ31N3lBQWFO
dN6nAmm0EQ3NSzA7455boa43WWu0s/MtAp2iwHKZt2rBUHDM68V0jf6j+B4woJizPP25oCEDM5uG
Q8HrItm6R9ZzbGYU0d28rusqKxlNLncuiTj5iP1Ecu8I/9MIr24Gn/rs0MZddkvPfUazmOfgK2oz
BzAxfI/LnnkCmY5VAmwpaiHS8xLeuveurj/MewvaW97PcBEEvF1esnIg5bpyupBpKrvZh7QYd8Jo
CeKtKPadZWL3LZiN81wCOJ0VPOuwL67LJ8hc+OdBadYMw9iWVsGWMcMl3/dKInfV+oqt6W8ffidy
hTw3OOxKUlRnkFSjJe/JN0/b7bE+EKP/O31sdCDzIYvHeaeSYbmp5hxjtZr19NLWD9Fzl2tTtviP
EbOXCP2KEONTDJblHbGyfq+oVj3R0qulyKx2MPC7/hN96jK4Nhz1qbbjndUSFOWYtUYHeqsLmXbL
VtfWVSqn15qJe7fLQ2qy2x0HkLW754jhD4Q+2eb/XnEmme7i/xDvDsDziiYQ8BFQQ/gMfGB/Hx91
5ofLI04fsgz6ff0cUYNKxM/1shWme5lr+tWPqt4dlSABytTlkHr9CuAz3Obnw9Vph+IaSvbLDBRY
bbO2HJeNXuRIPWhZKReoEHj3hQvZjwiq/XQp/5/mVfaScifMIt3qercJ9jAij7iBo/w3L1pzf3tM
+AGfSBQAgIG191vsLQhd4uQBgS4UGE/G+UX/OnIn+a+ebd0j8CDB718A/ja8RddfqeQUpC/5Lk2Q
z3SY/HKtlWb0B4I21+EJH03LqolCM9xZfvbbgeP7pLHtGjeWdWGPj4olFl8NvY2sL2qcHnCGefzE
EtEGw2f96l0e/wT/HqSOiBJIcjeVOkzqc47s38tcVjje1BS2fCUgdPlQz+H6DlclVj0EOC/N1+bn
PAZk5xEOr84Haorj/KhCYHhLn9+KRB4TRgjHZKZ/QBTAO6xQNgIaliLPf23LAYz4SpyBonAOs4Ze
VqpE+cxxD0aJ81qy9Ec/pTTqhpE5R2Bzkcke0fpNSzPdB8704UXO6lMeQjzdqaxi+2dsiamYl0Uz
wn1XcZk7kqnuvGsK+qjDlIQK4B/8VrQ6ZBRvdZqlQeifqj1uO/sxxds+SKIoZTYB+9B+7m1oZDUS
oOEBQumZi/r9n6JEBD6Pt/puWukFFQqiLilMn0NoOBOEKMwX10yl67yecqL3nF6OrUyGZE+soj1O
Tr4Bj3p+fSB3rIhiIoWQL3LrACu+KrsNNI0RUJa5k1lxMxy/7Ec+3WKVPIHQQEIBclmCUS0SFaV5
QSmlXXHRDYP9cZ9mWsy4IvNxI1xyNRwKXXo0KSGDE8xIj3195Khr8TKEXCnqQkTR+ExJBF4VHHLk
gOHmRuIgNq0XWD/GqCS17i4OTNQVgM++UOGOdcMfNZsK/jPcB43isu33Q937tPnKTg0K5OZhdiQX
3ef/d6gasZlURM9PgjnTDHOekkDnx7o6l4aTF0ghuDtPgfBrdl+tpWerrPVEEE8x/YFBp4r2l7n4
ZTm44N8evKuDucGzc6u4M10tw4ODSCh4VTai39OME7zXtmueq0xzjWoj73HAXE5KwA86ASRrhtmg
v+0WKRyYgSCxbk5x2elSU+hSH5/VoOHcTSU/VKHdg+l106NYn2+RzjM0pXS3cGVshS4FLVKlh2bK
kNlHzwBJ1pa2/vr3HKbFeT+UckkLJ0TI4d8+rOP/VIBGkayg4PWyuiApvFhNmN+Fev7hhsYI5msG
kdRmXXQeyYRrLH1ZNRCbXKqXO8Fae3yO0ikt2Gg8kBp2pbcmD85E9nehe+jeVf5o/De6K7sGZiSv
JkAoka5zIe13xrSWizQppepejQAvUHFtfO62GOI18Nkcf/GVZrHzQPK+GcZpafVvqaQKSw1KDL/+
c5rZ17oElwoPAQvg74mEczGnws6XJCnXhXFCAhozoEoIa1z6x4ty6U3spOgRWDEAKaZ0rdhA7/bo
ugZPMB/cPy37EXuwR7sPSIY/gRBZgZihM5XVcnM1NFSYB7i0tr8PL/UV/rJWuEnNpZ//SxkoYCpA
GJSd5ncSHxEOFdmRvHUkUnjplXB8dv6ymgY+LvZAp/fbnpKfWtqsPitzLpDveYL56L5nN9e7a3mP
Qmm4BleyrCEea6a8GcgLJLPm3fU2PkxM0Jy5X5eYQfOeon4sJR3xuSreVg9Hf/8jvW0kuUnc/yAF
sCqIjPbpKdo5IJ3prBYqfQmRmzXvYLauHFfRnr5/wfBEkftXROixWeCJhsvG8EXQk5gsDq2pCw+G
w3fOf20Nh07iCS2P4AhzzdoCyyNz9V7ugi+wAo7oiiRBXsDQ+3w9W2a9mi88Rpzlveb3yUtZWyyr
ipL1YwW+7f5L8LE7E5Tds1z3A3mdYFNW/E5B/8he7PZuM4HMsmlivVjTHYq8EQ+LqMNhIzMblasS
iCCFFiAgylie9F7iZDMWPuet4j4Ni3Ck7MkzoAckd47CXWPHgAgZRNLT5uZTABtUhp/So3iCUN6v
g+8vcWeDinplL7yhWG/mCYGgdP2QjLGGU5tccl/jUGwrccrIGEJd0edtLTu2L0dBjRVct7KwXTP5
LhrXUEiaqSM5NtAmWy1suBqlV2VuXMZkGXSS1KxcX3T8Vdco4DnZt46yRmi30l3++zi9KXFYEcl3
oM9VySj1EIaD/h6QLuSbOR0R6aLwwLsDAK1T1Ml1MS8YddnoVimkHqhjW21DXYTGEefGMjtvFnOg
YiKJEbrd5JLeEdcrwMSOQJbeWQ/mv8LuA+eiIkkK+vnWij6w+Nvw6LS1uG3DwYytsDgz1PUtha2u
EyZBvQexpm/MxY3rGyoeGlxSLQlBncecGsTn57H/sHj1UBBZTS7DDgPUwD9dO246/m42N4cg01E6
SBpEzf4OELDd2725d63RDMgWKvtpc3rpmFjIl5ATOsIegD0O8HkUm9zx/13aM8QjUzFwODYT3jI4
tI7NKDIg8XGPq0xa6tj2XvXYPya3RUM6R46hJuSQKFcj2xx5wX5YiRO6Xq8q2AU8VOQu8axAojmb
iYv7VsfXZ0qD1hadampTwtqVE05KgoU7g4T6ZQMKFJXYzFYoLyuHlk4U+v8wZolk2zTKZfhEIuKW
Z+x7Rn3xZQtzbFYoAzyl+T8wyJr9+AeAeMCq+/8zV0C2vwz1EkiIlDB/E065RU6N0lcsbGElkYoP
2Mp+2K8onLw+IoS5+504pzMbNptCChZFhjqzUhluLfAxzkYDYbkW9Ag829lYvELakCIowFd4+m0d
PmXVs0/RcG17KKopJGr70jwa063SwxUPdKRXwZBABYidFgEQuvBxYy9x/gSqnUk/jN/UdMfDa06m
cAq0djfImHnM8/UQIQOeiFzD6SHIZkEFdq7xXgUyrnoTarlSL8850hWoYICKaCiiQCmVFxiq5/br
7WWE5VkneYdmW66XgR1yC14e+xtEsGE/iwxzXTm2EdYl7VAf5gvJ6gqJmrQKqqTTjrHZSQhQgGVd
iF/SrcjZYgAWjhoBbMMuG/sGqZUEPjT8e21DNryFUa/KAKc4jlsQGOOgFgP+KvV7sXtWq48SUg+R
nmh5nIsdq1h5wZxgLO8ruDQ0HEMgQlC+AiHBDiskDuen0Wgk6Jp0gK93z0ruqAYOgtGYO+xT+cjg
nkckqjlSfeH4rSWUnUigJEm2ZWymREV7mxDv0CS8JhWqAYXqF7y+igbsfmMTb4P1Mltc9Ar6zTzw
18F0HED8O70Fms14iviYKv9kHoQm/ohz7G6SntVosEm9Q20zMjzz0QQlroA/FZ8S3wGrgkclEPyl
wkf0Hps3QKdnCjubxkU4E+FLSnDhPgqSiSswhBesOMPaA2o4acoVx4gwBGHFczQQpoJxFDtTN22H
FFm8eu3eOylmTSxpbcVfPOCFKd3oO0Z0PuE0vy5s87vkftn7xFKwsYNSPxNnDg3lTqAaCe724cAe
trygrnL5xYUECux282q0rDbhCyn0OnKfynZGPZXt/CZblbM5YMHSwSPFTb8ftA/x2xn8GB90bv3x
8XyqxevhIC7ikCAMavKKi59l1xcTSbKx7bkY5AAthO3VmzK3DI/VXvo9wnV5+LtDMKN4eH9U7blP
sV7l3FSpWxx/9AZoGRtVMObHXOSL4PZRNv3HR+de30/2tXBlSfIyj7N+AGEC6SiO5gFN0SxlrlYZ
a15OjBC9REsLs6Q2LC4te/Qzw3rhBqKPnodMBqoQn9iHF5BgjqqYSHPwHlUlHwW9jcykfxfUhkW5
XX8JR75q9rnuPPQLfVPGm0t2ujgLL3VGL3fhgNtPBRFExvmxUzSbylID69rkPj5MVuPIpvZd0Qny
RCdd2t4NTUbGe5c9c6Cgb9Kw+5FdyowXE02qCCHEcB2l9G3Q02H3uHdkjGxXqLqYYBbJ1kEvM/Hq
+KdUYbSyJRiLkgLxnAeRBprb6ekuDD1cs2UaNw7UWqUSEuq6muxM99oTcfeAEczc2TrhVMZ63E+s
itdy/0nw+OnBW6W9wxgEja7OdjNpCVw9gsonvEcGskTk/O74e2G9WKwUdaNy8tyEY+H28vZ7H935
zJDkXQrx52+YShd1VMGul5DWfRYmVXCGqj5pDOfFj5GoLlOTDAIN184M9oXEQGBx54wI/uw5+7gq
IqZqHW2p6r75cnDmE53h6xJDqTsnMUA86GtCW6JphzOzJwtJv8lpixYbgHlXeMfgZhV6Tlhm/8mh
96pv9k+cyDTCbguMhn3IxNK3qOTAgMeVhcFVWm6P+Ei9gOnGYrTa8w9wYrcpIs4dofZJvCrpRzan
er4ojpvusIzxNLlMpZoIt269Na97qpnMijqez+QTnQI2K9Jv2XdXw+pQaf+n/wqCnnuZCcBUWVFu
L5o4frW7mOZ1AHmRVI5qYD9kichNYU+sCOlfcgh/LvjqT0wRFKdBuuPo6y0IfHCFKUcWW+WaA3Xs
XXPM3mxJK6tyP+vkAsAiJtGY03ELR6fIleCKIyCc+J2SPB4SGaNQU/UhkBqK4inYgw4A2UDUm2R+
EC3O32a1Y9OJUeEAyS0Jptz2MJ61YG87EvWJgitmVC1Q8Yp9IsO6Vc8QxIeYGQDHiotFnNSXaHlT
f8EOvfooXFbe0ST2axNCUCtYE4qoGDu8rGnz/KbdrNynM+7WNaGF0EAzO/cEeFk2APFEgO9+vBnO
aIi0rM3oN1IophaKkdogfbSHU7wl4cwO3+oq4i8eSWzwifFIp22FAUHYAv2azG3G3kRpDwG6u3BI
d0EduR5MLXngG9p6EyqCd3gSpFXnEhNsbfBSrZqWwm6tS3goxWN/ZbvTMxknKAAAt4O5Tmt+xxl8
+vPlDfqQ6Pymy+vmusuXX5I6VqCWrbfrKptIoIy7j9Q6C8yr2L5okl5786tZ4e+dC5AAOqNn5/yH
K7kvaSwv4f52w2msXavGGRmt61cEAdGNctQxHq/tEh+YJtQNjTmqisM+0MbLX6K+FiQrH44iGlQh
rBfWqs0iouVg2rvBBBP1YleuxG4rTt8EGZg8sdUUXUlUkw+HQAsC6giYTcSL4yoDvmVZtqg7WA3q
Chd2Jhk09o2x7RMa+YDgZ8PnAHT44yLkYek7ToM2WT39X3Og0ff2Zsm6Gst5YXbiGvZvnUpO5571
kzliLkR5NsuHyOa8dXYaig/IS2d51Ciw1p3j6mU8vVyfcBTvX57iKObTwy1w1pjmmUwYPwGGftmS
KxnJnFv8pkRSAeeNSNwN1z0PFA0LqJB9Pp1sctMsRcQwAFR4hPbf8JsLcLNXlFa345qPnBeg53xb
ZyEnecHQ3MyTnQy6bZ1y6fhcv9nNJJ9Ayt7Bei055OUcMfxsMJ93Blq9horktE9qCaux0PAOBe0u
BMGkKmvbVptZFks5byMToC9YnJ1iiL5u7vuJOz+3SCMu8iylgn6faxKxTqRk9jz8OkXyOtrKIJDH
npnkYJJ7XnzhzlFwBET5BmQnwBGc7F3f+AZE7QUQ3bEe5a2KD0fJNbYzKfT0SZEkbhB/rbZo7ka6
9YwGRNRERdsdYNDLHPkRYcwctwvG64QqdVv0C1hy5kIu4vNhcJtGehHn+uT0r9pb1ZbV2iNU1ojR
syrq7+B8a4bKCOiueyLDWRnpwuN9buVE8xvIinSPnU4a7VW4oFE1I6mwk9y/ZgP5lQp3HSF4vDkV
LViEvnGpZk1/h/bpCHip29FWvXs0vbkHHym+Nkyc9686RVR2s1jAV/xpS/+v5GvbiE6dkgCrKX2o
9yuc4B3+Ge6pIJO/7ZuAw5D1F4JQVlejJsGFK9muv5l9gwl5GOGzHyJNJPdikna+2JTzstXKhKHC
JnnFG/45ZW+jajSaxb9qVP3MtM4Y482CMew76BeEdstg1Ik2RdcluaRDpKmTPy0LMKiRe+Q4y5MA
wx3mMPJ3N3nzsnjX1K5X9iSUf+g2rEGOh14mzP+mxyXvy8cokUdKh5EPaFLOkjARMCWxtSJSNvPP
2JTbpJh0a65Yx/wV87X7T8C/pbgZFrg8vKqpe6WNgZ2pCbb0+EtptPhs4DOhg+Oo3zhFBk9K5YIq
j6o3KXuCMtNHkw7YX7tQ3TxnbXFGVr5j/M++eLdCM11raihvfAqg5Z4KyEZv7Yh+HlH276laDybG
owJEwl91E87hrUx8/cBOwX8nVy5DiK/KPZlRMBuK87EYw7vQfGlg0K3TDJxO739/s2RVXU7+4NFV
+hYGKxe2navUpMmL6jsA1ahw2GSsSEnlzz/YrLuz5hQamW2wxz2vBCtpwAa4OjTxeX2JmYA5+IUV
Jc3w15/2B71W9PjnIgTlYMZ6VqKEupVL4Tqyqz5x5P4DwxS+RgARg8D8XLE+h3TqvqrFkuFuBMVk
oqt2ve2PxR2IvO2Of4GlE5txEQPA9p8P83pV6t+7eKtWa9Mn+FKxHQxGlplaUZpUij0bF7Pb8nrb
n2CmJ7D0+7ARvEguUBMgz3BXUli43FvCoIMmyp5X7eNKDc6woVJ9gZlrvk1TDDEeHIEpAc5GiIkC
1tPGHGkRlgYdo5LPvbIYjt0GNPfRfQX1C5j8g/ZbOn8T33ESZpZHxjNE39WQ9yN24Tl0fVq8kL6A
V16Hs9GaQZKtv4nHRyU0pDIQhWOPheNeNwm3ytF7f65aqyiCdINH/RWrl1dMGrYX2RSfNqMFC97o
gpb1xxWY8foAohF6kQgRAbX5kNZ8epASJeLhYNpCsSTgkjLbppECT4mmp7FyOtU4Wa2V7IDIkfGG
LI68LpJEZRNXxbXiGyTXl5zbA5BuCROdkYgd0kN9HLFdLZ/16s3b51uCxdORUV6k7hIBnji3tm90
XRDZI1isGuruZAfUb7QkIYaLQiKkasajZWoDNveLiL6DezfgUfF7nefIDYdW7l/tB01kItTYoRBo
oO6NtggLJHw+y3yZomnJrnbizLotLkt6CLBF29LXm0QHdBdt97RYmLw1kjpWnPd9of62fsYCKcdl
zzQzs43wRWhWg/y8eArTZaG87byDGNNkyD0oqy0MObkcyb4/Ka/V5UWMiRqbZGpsR1JxB3R43Pf1
Ab6DVFHMiFmUnBoAq/q1iZgxMKtCFYDb+4b2jAjMakUUFow0wqmKacfEyya0KHZWIU110c0SaE7J
cMq2HQQHiTmtM2OzfpnIw9vCPTXFHvvwC5PU9r09IGpZfav9mc4SympcGk/ZN6Fgla3D/Z7ZNwgJ
kbN+whTG+4mqGrfaQMEB9BrtC4H5FZch2iCcTG1q9r/z9mYtFHNaUmKb/g/Mvli0HuYM+j/YSv/D
QFLtO8EGIUNAovVC3cpfcG8lWeLXOuttLO5OgB24aFsCOGxlprqNAco8dcGcgXh/ql1jwpXCNzuH
MHWlzrW4EhIAhyWAOTu83gjG71nxnqV2+zRm+lHS4PnfxzFiwo2qKrMQrfaJ3llhYpVN5FjlIKPz
S1I1MGttleB7gg93hjFIvhcus8VoyV6rZrnk78128wqbTZ4OTpUHPO7HnRk9qFyUQY+ZXUoYQsvB
NDhX6s44ybHvim3XUiCM3/00OPtCF5P9sIaUlBfBJEhQMMSiDc2Jru/rr+ivxeo/GTI/KAppKicj
IQfAMLZvKm0CEMnrWi6T7PKwK6akfnPxm5NYvTHNHH2ONB51xTUkQcJP3+5ayfmevaJHvdnOqSBS
hUiyA9STbvNG3HWOb3ShbDsHvCOd3w3g7aUbBeA5WSynv7rbI6ndUmHP3xwnmXyD03SbRoXiUMfA
QA70VlFsqJn6IogaG2uPT9eIht9qogGIV4yP5nGBOueZP4nKDJys6MChEbGAQGMXDVgazzSZQCv5
pYp/mv+uqwOIJnjfs+FOl1Vj8YDn6NNEHTiBIpkHjf/t11KYBV8UKuaXtQaQhsBLLJYEkG4tsM3x
p7/Ht7ppVlpnPryykyR+sd4UAIukAbcavI4DfBjP3Szy/UD880r9C9+uG+Ct3Y8w/t4EC8klLZTY
jvHJYh9cWzyjnTjcP0FiYb/6Yr49hDlWCKdYHdWqmGnHB24qYtn2KMYfam/KpWSOCIatEMxK3HG0
jshsswtwgTf1pBldntxYZ5oEorrpkCKxph23VMs5k0rTWttmcBJwzagW1z22anC0DkleCKn8eI0v
yaOxGkVT2tw3AnUBh73vzZgJHYpr8krWuJeHdoE8Bv7kdrbG0vDO5NRFxqp5pWHs9tQTpdd41O3L
uYdEJXEE29N8g2MSmW5mAwdqu0XAPOP0Mj7Zaw4fhcb9mQVxx0TT7naQcIs5YzwFtvTyMr5havME
/H2tAZriLCDkvJadaVZ7wRPzmhaL+MUVzSpIxkGp/8MiZfEjiozOk7N+GBbVg3oHsmbJEZcJVnto
daeSW3YurBqafPfStvVFihVicGAhu+bwg/HaSMbqdYg2etMR0Cm7TiJtG0bvb8bposjLW0quiE8R
XkGoznQz1+3hV37RtpnHXPvJM7eanZG1JpLLpUlnvhP9QKuIMXJfYz4vO/UH39wFZVCy5qIG65jM
8AIVRIikKN6uHOc8EdISOKVTZOI1Z2NDOSgc5kGdD44R1DoKprzniXJym9ZWnZQYFUcUHbBHI2en
+vFhWa6SP1QdKL8u1NbboBg6LnX0BmDRe9Y/H5vYhbBs++isvVJoSd1/WDik40pba+tJhH8SfJUm
Zq2wiMgOuoKyJg3gnkSRqmxMucGSnKLiSzq3aV8PPfmX+UpRvo1Up04v0V65K1gc3ETn5A7Y18dJ
I1ylE9KyA6Mdc01bcTi70fes6JBH+tnZ28P7OpDjnv5bO6fEfZbDr8i94LhJ/aAxDBUimgSEK6zy
F6cDPF+tOrZWeQeospqfCjZArIfFzGXu8woZaOL4vazSyAcxylOX2cL27ESI/K6H8EyqxSKdZ92f
9uNYpMl1BQSR/faQ27X38irQrj49n1tvntFRK9QAqd1D83zEV9mbH0S57qpMnaF1+pPxd70etgIZ
GraJjaPptYOz7E9j9tZ7PRnqoSul1bev7/xpK0d1QMogf3M0nMt//sZr/klujPzsTjuNp8heuiHO
+gz4nYzikTvipHCXuoBxaWPWdntDaAkbHMHBqhE72TKB7im6zdXNYq19IFcX9RxoxCQFGwubCkXk
M4s6kCRG8SdRnes2qduOOGWad6f9e5PyJIqAbeMJRJEFUCELyceHS+dhQWXSqigl6rMvGPuIiagl
JG/qVGEFFCgMdaBIzvHVJRb6P0qZWVw+8K3nfZHzvWITuUa/La2K0curGUvr/TxjSyMNU5HGo/5f
0JYbGGcGFrkHPOYyzTZaqK5rUoJxc9n9gqTgiylaAeunnxQ2RV7viXn9gZvU+SnyEKeALsSrkeml
blEZE6BMYefHARbdCXg9MQ4SdvKZhU9zD2A7o5QKpVVgnhvx4sn6FBG5qBbQOwoNF1Jtm522LX4h
bYP7TPg5rhp4hfKcUnqjkDm/7avJ+cJ4iAYN4HFOpQPAgdvNaRSXCuDTJfkQCOeJwW/i3N4RYcUN
u7+vE6kz3yjheNZi0rpSU+kqqmHqTDymLOvdUmavJWXGljM1zMvcipnyEVrH6HtZFvZLclW+w1KY
jukSd9p0Loqfm03Xd2oUP9NNpOWTOvjRcVn/9xnM79hSrdLbRdBEO4GSc8iK5/e4C7YDEdQecSAi
EA+88dr5v0lQ36M0/fp3ZNjhPT6pwRsBEU+o9KBVzAMog8lkCiZknKNu2iQQjfhPBxGNszD5MuIP
M0drNT4zcSaYLAd3Zh1mD4B8Fjv6KaKonuCAsNDd+7dT/rwKODmjQMdCbPOaRCtwYLgW6ZyvSR1+
9N8Gl2LfhJr5+BfZpJbHC3f1nrKC1io/TD+fzfyM9rLLL8AdZRV/2WmgcJiUOdXfCtNvQ1WD65GH
V2H6kBqyCOyrrulAiPRI4PcJ1gZg7OEEVEWV51OhRDhUJFBvGaQhP26doRNefi7ZVfp6wWm7CMQU
xVfPeAraZK/PgrLiAOx5NfvIm65X+OZEJ8bOYsQYRdiElf5D85t22kmNxhhDULyjG0dX/6BJ9xad
b2XP68CL9uIcZ1ivQwOhXIeo5/GNKAooL4vEYG8f3NxDDpgDK/mzGa+b3vR92VILEWsj25Hj+TXu
h0MUDmIIO8Ml09+KRqq+4r29MFVgHt4AXUnceVT+4E2bW/VwDdoyS5etuPDVoWWeFQkHHY8qSOgm
P7YJmlzdPQO2sNAAFKD+PYWBaXEb9hNbDqkFzNZiyjSHvavOhLm44HYntlFO0aaUiDrfu17fk8cn
m5y4A8ZrUWI22lUe2ElEPQJaSdF+L6iL39DNeCWJWHCDEwOzYvju9afLsgb+ontRDkvkMPiICkhL
BHQFas1a6jSKjI6jpydYrvJ4QABXYob4nM3ubx8skLeBmr2G6B2C2uJ9p5dxFrRcrAhs6nzLqVVw
T5DMdG5Xdr0XJ6NOxos+YMjetbLafj6wJvj8HpOmgWUvvV6emEbsFcqHTsQAvojdYHSNxMuloDx+
4kFOiJRnD4ikmfRmyhxLzy7hgCvNYpIqiymUV4HvlFC8TjTVgGwQtcyzSHRdUw21FBmQ/33ztp8m
h8PrIFYT2CW6EY56lt/VqodJ+IfVfPJtbXC2aV6Pn8RiDVSkeQU3I6m8IhaTo5noIJAMqNCzD7zL
+nj2hn1uZDHZqIQxDgCck2MXLYN9mYWOlT5diJpRFm4e3eNdRr0Ir7W7Rp7xwmsaIoaLrkhmOdfr
1q5ATVYT8x21IZuXyltCdkb+nPNJqwFpUOoYtmfHyCCfSuapZWSinD0m9jzHGztGvgoSCLFZhPWX
y3YClJXB6vI8t5EO6ZXPU43pNgVVQOh/yF9FkdMzSP6DRQujeyjJO+vcPhbR/t9WVZEIbvcPasiY
BSMo9I+edA8YWLFqYf0DBicX/ouhZBejlkeqb1UTzKnqDkVFdll0l29vpH3vp6JlDEBEJvpV5VzQ
3A3SbNIxWsFr4gaavGlWmwnQx6H0Rnh2mt32ixHkL5/pECKJAJ+NVbLVbOBYF6VJq52U4rAmNYEn
1LdpB0fDzhuOltOv7u14btaBZMRWYT2wzr2z7L/JmiLK6amBGY1cFi9tb+IJwhK0FQLvoBki7aq5
jFAgW0RIkFt60aT4Z1FaOxCc1PTdp70qNJeO24a6mPGBFU4gaMcaW/zIrtUp54H6OiDZy24jTHIN
bfallmP7wa3ILZI1UCGWzk7R2ogfVR4YvP0IKsxcv5r+EdomppTIBiWJnxd9pU0z8jqkds+dvfY8
Ht5wJ+dHOT1Ta8bX37EtFnF7157f2HCC2mOYdPKG0CZijHwUWkunLCFUdRWUC59Fu/ZIZRasJSyG
gMwSCcca+C1Vxtq0C6bGp2shvysNYd7OjLmFSUdpttEMHRwcNRfADv5ls4mSpuJ4w/D5JslrtgNF
NfNqbTNiBPC/MMK29vJk7RJLnz+7X68CXk3FSFLRnLy/14YYn2bqI0C+RurxqGVCefK2DjAv83/u
1cdmo9Uoi/d3Ktj7nGhdgL7Je95pWFf18GxPv8YuXkZw12DQSzk0hJCO40JCyrAtIgYgkjfKUPD0
etCXursWgT/YgH5RBIMAEScK5Gxuea3kpv8Pm9jq/n0vOvmszSdRBhDSLOZ0fliJg3rEwD3ETtpE
4oKKUEf1hxLfYTWdjbSunGDjKuxhyxnrW/7ZHqdEArNVX/Iry0HWIbJT0AGfAPM7qM3vYbaWDf6r
dcRZs/j0VDDaib04FyKdXlDGjgGC1xicZLKQHF0w/48rgZ4ISka4U5M5ilww2+tbZg48kadyxzXp
tunYxrJPUiRyY6M95J9vg2hxjSSc7idECGKjaMej3AIRpUwPiHkxiNpHGIUcb78DLKyfg+UMqYx8
cb42k0K8Mly7OQMgkE3Gof6ItzR5xJ7O+sWIv0mR2ao9leMPlyanM98fwjBm2vn+jdFgDcM8Z/aj
WN290oY57ZwuOeJwsl5dWMskMYlkmZUi9OjicnnnOjE5s9ZObD141m66UrhhjLdy38TUuUP6vKmr
i/ezt/JsKccpsDBVk9+3FvrKkCBvOpNtq1BlZlyB2XFnVE+X6yZ/vnP+IZodqv37JyRtbWz2xV6C
LC7CN86E+J+Z5K59Jds5ZZhHan65W+IwEDFymYDzSI3ZHmXGqAXA9Xd8uLnjuvTuhxd0fYehfeSe
IipVzbSp2WewJKemtxwkt9Ql5Vg1YL1TQ7SoMKRnmiE2Wp9VrJlQukdI+AnLZF3Td3UX/vYzS/HR
6smCI06vfWra40TO3DuQuuT3PP0VZF7ILdomGATPRMpNjBeC4nlARLAymWh4FNM0Y9QOGa+n6BCP
tcrwdkiAVH+muCUIg0kg8x/3lTAH4T1+E8a9tV3YdCBk65sN3oC1pgUsQLko4wCtyNkgMd0L6ZAf
fipoqFElLQ8oHYAPQBk43ibKSMuBLBMzTMFWACdHPfhacmdqkhue1vstxNWP78tbhesrrsV+K/Sk
RT01l7pd4dmytVBq5ym/aLNHrlGG33Om7lGaWFXipeX+MCEtrUVcWY9Ch1GBh4wVLccVJzNIH+Y9
MrS1mY3siu4IEaUqs9D8DgI2HU4TT9A0pxMAKpWYt1MX6Ovwi2sdmZiz/LzsQQt2LayQUAeT+J7u
Oy6+7/H7JWZP30WFbCzk5hlemcS3f7G4CiMMKwXHFWySi6l+WWv3zeyTzjzLXBZLT4NUU3JV1D7q
mXu2L2J6iGVEgjtHqUGYrRSIgiPoPvyOtlDsQpj4/WV/bAkhP94hLVfT+kD34WKR3yVOsB4DGcsa
x/IRmiNXSFSxYNNOrd72iJb2rsIjSlwEJQ7YjpUWSnm/41Y2Xc69+lQRmJGm94Bz7LJGPucTixkK
ToMDjgYdM010XG25P4jF8VByxR1EOW9PiV5NB9bVc22yjFyc3xhMLpTwRPcY5ZOKiL7IyrYxL8mN
yjGtsvgK7HV10NQzV60xlz2ohJncUxwjAkUV3Ul5ezbnuKCWgbvMXAgvi5Dwoh/h1SNQZaCVBNVv
cJVlRGKBSj0G1o5H1KxW3FwhP/bBYkdYPTCVuwhdVnTelpPh5zfOb912cHDcLgQeb1lrB2ISrkHN
PBKSGcNTRUesQzElArinWoIa7mIs0MJzNKtF0svpz6i8MB2oOictEdxfarLa1IDlXN3LYcfOvwuw
odkcUvuRT1mNgUXLpX8GWccWvdx27mx7r0N1rsjyDOt1QO7PaQQsiNB8v4TbVqZALLnTINedphRW
aDsZWxYpuLvbx/E5y8in0S6XWNu/cqVqG9XCJahdEnVcdiG+fLw+8zqxlS7w7fwxszl9PbmCCtwO
RRLOPfv6rETpJop3wBQMWXuTs0pNE41TujuisgJaoFaftVBPxpkGqwhOZgP6rg574t98posLTTmx
HPZ1m3MH/GkO1La7w1CSESalVCxI/3LLo58Wt+Ft7osYWM59knr0h7jYh7XyMTFVFwn6pI0s13xp
CFNH6SsR8hmz1BVwJDJh/UgDXXDnnX9B5fzJpJmDMn9zsjPQ8j73pyTg0/EOUuu7prhl2jT5n7oR
ovjxfsF4E2gs3bZJQIIgZ7i1bVUt0C4K/qre6oAyMDdGRdEj9Zi0Z10e9SWsLPOCC79VIWo1mC16
L5PTWgOqGbeGckZ9yjiAj1ZYZlOPePtnYlUR1lNi2I8bXT5Up1ga0FNecLCq39RbgHUVaGjWyPtT
YIMhiWiZWUo3uJZ+XMc7KBL7fLZuwIEETujKUNgtr8NXOQiHySCMa/OzKA9l4w+2+/SliQabzQy9
D64D9fKzOpBGaQJaEj9EZlSL6NJ3WY7vSvcAIMlMdA4FQhIi9HUmgmscN9N2KioZjX3MwfY8vnm1
x1TWfL6MbPxUGU5zkycSarK6pQK6yc+hJlEt6ZOLEYKauj61H2wIGO+MzSPkag63d2F4KgTEjyJ4
zXdbedYHl1v0FWeSny9ZYijyK8+uxKJC2giP2amD0plu2/suBCva2MRdU66tXQXdRRVMW9zgwBIs
ZweTKoOKcCIs2DA7rtvpITOjoow2YUE7r+IMxfyFW/BEnGoHmgXI5YxSBwFxbr9bmmMyqq1kdIVk
sWKqotKuDdXrjecvkEutTinyV12SmEThh9zbQPZbTXJJ9Qza421YvgNd2bCyWpSnarYopTdkBlo6
W0VosMt+/GwQAJouIaXEkA4+6/1eyZZR2wMpvHHlvMM2Orvspn2i1A0tPCQe29bElJltc/vnTEWD
Qg62YGzzyTcfHaEN5Jffr1tMdpCXhTzh1M0xibsLbjvjCRqOjEb8GnEY2PlLbYD+2m30DF5iHzzx
rcOiXEb4nqBFCGKzgg42Zv56m2gTP/jDX7EJGS5DZ44Vt5kLiqij0l5lvsWz7IFX+Y9wNzrMcDjn
nZYMhQMFMgVTaSBdm+/h8mLB4kUFXrXITcKW26pyVlCIU+WQCOweETciqueNLqloSYlnn6DSmTN9
S4Driinb1LnTh0StLfuGlpRC5FMiAIK/Wz8pnhiUB/ZSSQsoVd1uJV/tH1OntIV1K79hNbd1mTiI
AzTwFhCIeSzZ6tThF5tj3Se+jyiZ7ukO3G65w48fRwOWKNe/9ckgwaKKdQW/aPkal6PbgsQpIx99
C39oTj8Cn9jiZkY7kMuECa/6Nq4slCjF5/pFC+8helO+KW1KB7ImLbRpZIPNUE7iD2HvtWxcPvAZ
/mIZGSSKA69YkkJ11Qsu2CliefbG1/HGtKBhSPyo+Q1l+AmugoyMY85oczm4jiAZpthHU9jcVPBZ
dnpxYfEWDFkZmIZcC3/LI8KnUM7JdhWaXwNPba1vSFJBGNAHdmitRIRFySKfnud/RMnP6K5Aa1z7
KPyIDB5tNCllW6OjR55s9Mr6lNTnUt63cYgrn8vpP8jDdDniUkCzOw8Ey37x7j6RWtZ1nxX47vd3
gNw92imqGmhYhIM9fO4xZm7SZNwoCwR0c7q9YGAG69iO9FuhhUVGV64zaLFflGUUhAAd10yzTv62
0oNw7YB9aOyYwnjIdGuAtTF3e+a1a+nPnZ/sRxWcdMldh/qi5TiRCFxGmzWXTJcyTAHu0Q/xakZa
3A0/zg07E4sNrXwGNaBuN+9lqZLoLORUtZllcbxgAxKL9XXcSRDET4hpujbvlFCDuZ7vET3K7y/b
2TVuLsWVm3xZKxRy4bGiF+gOqMtFijVI1kU8i/DA9ciGMX4T2fViDVOqWgwiTMYIzZw7Bf2V9k+I
iiSNLrtYLwXPR9JKTuER4QTVd5EXC3wyy2EAby59ByaNgLB5AKXAF+hU8+0ml9YNJztKrmOcDgXE
+2ZgIqlr6T74oEvqXaO0wjU47A9/xDrrb7dYg0TolMiMbxcqBM5XeC4Gwv8mG5eqN6ApwxRpFFDu
hh66xVWMM+uZAzTKuPRSmU6Ytu2MCv6TJ1D3KzCSsStUGzz8EdBtqQDm/cx+uP9kzsC25qWS8XoG
Nx4katTZSoiOGEl0bK91DZZNWURGzVn+yKlCyLoA4noS5tGQctyRKJ++lHhZakMYkmHTzSeGCMvC
0Clz6YUqi0d1tkghviag9UvGNH84qHaMTAGUhV7nMVS8SxJfDfI6ZWnZYyL893fZHqcZPoQS0pcH
o32V3gJejbIS9shr6mdyyVP07RsAfmdTeE2KG08x+spEJDP4dlEKvrUHgMR9rJS5MQWpIhGeCcE2
VwXlR6HpB9nG8XTxvu+WTXgSZSMA50PfXpXBawV8/oQDQ1c+qj//LoEuULMpeZ21MHWgD0vpFLsI
QoD8AFtiH0BgfPId3Ts/BkrWWisz8e5defit8xY0O520jzrhcdiBy58Grd4PzgmZjyUgCx7BFbbg
O3i/5cenCbjytIqdmAdvMZ/C2RQxRVhCuVyVocN8ImIQp/2/UD1H+IAwVhYHsOwSvE7ke0bVWcHL
NCxTlL+BSdwKbCD/+zWZ7ezgs7QWu9Q8eTFvK4IQFgRIASlwbF5k5UPHOCvzLRgXGSio5eY/0AY2
B3sLyxhdmpz1PjrSIDrovGyPNo8XUf+yVOdA8tMCVATvw09KoJwpA2JBqASsp0t4WjulJV117DNP
rwZ8I8fJyvoas0hvRZ1x/QzfWBXsMFKN2ZH31fZAGAdm5wtytKjmEBYV5TVugDeoYWZCv8RJ7cHV
GV+q+gqsqn5QvUOYMAzPft8UCjSqvTNkl3pWKh92KG4P7bYwQRhYmXtje7X74eoge3uzrTL66b2N
tuG0TEclE87ELHpyMcqOUYmi0m4IW/Mu5nEJ0du+SOUlCCMKKmmLLLiOfhRe4brAn9oI7ZeFJYAU
KhoOCUmPkufsCQDBZWiXN+/6NUgreF80eOulAvAsD+shgrEuKQG2KF7mZutuLrHdEa2lqtYJLkj7
n8mDakqwSImTj3Caz3XE3US3DZajJCE8cJoN3t/yZIqN7F+8G+udmpCsJR+OtX7yBugmHz9Yx+xo
XvaJF1jWVsUwh38+lapFsgODjboB1sy2yCgn/BBH6LQqpUzHObW0Ur6dM3O9tJY3mB0KW09aDAd8
fxO3nV6vwI35ipF/Liph3m0AxOUfkUoVsaKMBNOhm0/CV4SSu/W8kIOLc2bzEgGSAAOejp/Susrv
XBD47u8yNDCTlmtsbkvhVOz9pDpbllREq5psedQKdFp+FRoEnV2JDx4MyJGiart+4Zy+NWOCtZCw
RKsM3rOBKbOVD0fgV0AE++ukbGnxO3cCwvef824R4FW/stzZEAXpQHVT6Es2xFuS1qac7NNBtGDX
1jvEDfyJ1ezz6Pvpo04jXniGJ7fTOw8W37QX1FpD8+4QYtIdHuvhWd7HX7gbQYf7rx/WTgrhpSpa
4U4vADXpAp5fA1l//ZS1Aaw0+obzDXPBzR55K0osxw+elDX2VHkYw8NI1wlljvoBSB71XDOUPdcD
OD2Irz2jNPUDbd/oQfL7GvlFd2BwD+wQkWItXwr2tzHcazd6isjQtxm6qqaoSYDql0D5F8CADsql
vUoR4sz5+mZ5Tn9vbMDptOUBkV+Z8t39LjVuCJyrnzFB1EP6I4V1gscEjvq1ss5xMrYgobpFedxx
kOWuRVEVDwQxu3i6PWQvMX/JsBosKjXftE1mn/51R1njBtUFhQ4fv1Wc9DvZ1LNMrMx45QMAFXvD
B/RE4dN2revM61yqx+VwXqRm+bF9yyLk0jzFoI7mh+h4weEMXSiuCkpjwgTP6KnGXFl5LR3Er28L
bjGVwDiW9Z5cGnTldsKiOLLPsrhQ5nUppxF2uJMBqcsJZd8roHxue7ygJZAGiDG2MGL1cb2LHg5i
CO3fbBNltJLDkmHjKoTE/A9IKl3jj6WqkdwjZKtn/wX6AX9YwDU8li7nTRi7CJVjQG4OauVxSuT+
yq6mgorun1D3FCs6EBUS4PeN3kw6xjP69OIci/cLOx6BKZX5uroGqO4SzdY9w0G6jtrXQ+mw/KIS
1jCxX1cf3wNj8i65YihslwP7L3So3491vw5sWV8BmKOmtzeYkJDdpscOZRe878WfmkLW38YRanVD
ar/SW4pwXrrNbRZEsJcmxC/Jh13ntg2t2Ym6rtywsYddeabSthXZY6uZ2zqWGavAHMAo7ItugatU
yBwlXEl71z6owxrWBsrD8G9eekvgQP9Y4v3I7G6toV2dQJ6bRCIwwNZfv0gFAdAl+vfhrWZtLgt6
Jhp72diejTr3XBHkp1wamP9HsH0ZIozE4zuaEiXpiNIMUZ9q53mNxQKPouE/FRymYADBQ/J0+Ngi
LBBay2YdSCA1CBT3CbwKtYqZD8lrMM1W2AJ7FuDCSCmxAJk3U8dkFu5F66BFsbvVNjmi8sbxefj7
Wkmee7vucoCZxJfG+KW4Qgdx2kUtARYZoXsFSOrvj5LV6VBYh0pV1LRDy5fgiNzC0zdvOW6JM7CB
Mfl39/k9ktWXB4f1n7bfbAhtGzxcv21BzZ0P3KitHK9qW07taqV06cBKOpL0O4uzzYagnDXLN5ph
nLEGexyT+Bkq2WuuLwqzC64Vu0C9+KclRijZCB1erzUuZB/G6OYTQc93ORgQynp41jR9df6QHTej
f3aQVfiV2H+EZikaP0oKzEbpQ8GsnpLyHOBRQXQhMlvG5lhpgYrOHWWw09A71hYMfqIHjLxCeCTl
hewUVGp6IXV9SaC+t/h8foB/I5y1FRJbrlc+lxfG7uTKwrUrTE/9jASPzDyPfcfzBKZONN8enJub
8rExmvYnBF4QUoJWGNMBWYi6QG9XvZ9cgpb/h96eOPBVRC7ZSXihsHoBZNXovFCkiPMpqWT1k2kc
bQOpJgXT8BqxRuYCq6KV9RmnVYduXe6xIROc8wq9JXUvoixQJ778brg2oLKlPu46n/t2Oeix/77U
m2l6jXKCaF7gYg84zozHDJfQgiQHnc0c4jHNnQ7mhU2i+zOAxwtcR7MS+QnjdaMfVYHHW9N57Q3+
wICNZdWwchp6nmtAgdrjYub/r9EnR5RT7SFj8h2mLWBOnbHT3ARP2zCZYTgYzn1W2rIWlQ2PDkQd
m3TFAY6MlQtWCXjaAcp/YsOpIaoC5hnMx37kQhVG55Bz5cUr9RxSVgH62iexuEFOGdcYm69OhqXT
Rzh2+JcsCLVDPe/DuJw1ATH/zvq+pBpRNi/eZVORg/xV0iKOC7Ltirtrw49ujBd52aCHk3u8d236
mey6Uqc+g8kUPJ8nABBkh/0tAcsQVVOZ9fRSiURckSDM08y/+MikOsvb5icTpzPPb/mC0ZItZ/zd
htva5xHGIa37pItfcgxC4IG+3aVVfmcoEeE2C6VaZMMSBaeehUwS2++ZZ+VCUgQPCjmkFAyEY9c+
fWJ0uZanOAZ5LNF0ZkFsA9ITTQtPG3zOD0ZVWByLKsnudiTaC9gGePhAYjyNTcmqs7KWIt3IGYIv
Zj/espuM/TLLnJUzrSjO6IUXr7hfcN9l/AYPE4JoAnev78ZQP8kB42CCOZL2lSRgVi+yT4b2vMc3
pgmFkEY08ATpkj1vMobhdMNokf7dNGmNhpWPIgyJDoFxty3asqGkRXBCTJ3zC1daAyLlUEC0SmC8
W6ghXv46WpPP3dGQe4q2yrfGi/O9dRXWCYFB4wKHHHV/5cSMtPpVIZvkD5kZv6c2Q3oBhF4cab2m
tcm5P+rIpEp4gE+eVMqKz7NNADIj8Um/N3scr5JGsWBkyz//LjSrLEXpzkzDNyQjPVVMyGlWsQ7+
wqzgO32/D37JL0hCPx+uuT4BoUJr9kkZmNwo3TJaizTccc0anZxPStcq9eCnjXSHf2azTRgmYiA1
w9x1oPcyUA6l7pyvrO8CmAPRxHAxhqtqidOTT0g3F0C9TMza3Q1C+Gej0NTlsK6uoXxb5nIxPggL
6c1E8YyrS07TTSxK/Sb48y+8zrrsuB8LiRw4J6BkMFfYbDd7OGlNfS7UTNngoy+WamsrF0cy0mab
w4aQ5PTN7HfdrVcNXk/iY5IvzSdmc7l2bCH15CxowvEaoFyDRN3500Dz2S+1IB/0ZUT2CWZZBdGL
8kc5FfiIw0z7a1LsnBtXY8DVzkgMqeMviGsrR/UURsxqrXhygyuRWHyS8LuwTA2/8H9ekjs2Pexh
tBCZCWDXP9e3dn/XK2hEMzdHoyAZ/rSUDIXT4TH9vyjR+bopSLd8kXXiFXA+5xOfNpzyDpbi95Qw
WDhwq1lrK9j4b0WBE3iqDQMTPk1pUBNN3Mg8ubiYMZ0QCv++GByz8FTHODpDoPQI7cC5G1cn9yUD
cltV2m4TXWhM6/1HI3U87SRPhrgIo+xwrPpLm8dRX8nPD5fc43sam2jSCc5g/TavndLescCuXQgJ
NDF8x5YUMBLjmOCeUZLK0MY8KFZxk2QzbYlztRDWtIYdM8Uv2MF4oH/pTbpeZtLYmLxYUrWrQsmS
0IbK3Y1owhgXMPKdJwBcYssYWG/VCJg+K8JQdzvK+46EJgGrTYdnds30LgEBVcurTIdcvdfUTO6e
Da3eJm/7wp05nAZvPXi+JYucbHU0of/Yfj3PUDOqsFqXlHGOsnxNFlGIq9PZa/5IsowonOiCbxzs
fVutEbArRWIC5ZRXkJjx6pgo+lQYlxquWQUVWw+WUeeU9WAjEmUCsQlIFwqdKkz/kZUit8N8W1nX
S5iIa1ltf1ikNi+cn5z09ekpX2/wWi1ibaoLljnO3KlSbKKdXNxcyO7wrumwSBRky3N/N2mmUsu6
tA2umxtEq7WuSpSLl30VxcV1VUNM1DpD9vqtBW4RSv6G4ZAnVj5Is6DDzITK0133G0e32I5MIwr+
rCbLiY2ZnRTPJ/aiF4cclNGduMl47kZD4byREjCmlPs4iIAtEnKEA7Fy9duyH8gryKPUqFpe12wv
ER+QDUXKrADsb9RG2cBRTOenRBCLzDiQk9H8Hqel0rB1JY68jA2GzFL/lWUlK5Om1OxhLg6fbxrG
01IIMNn5gsX3pz+Hu4Sloy3uJzEJkUZq9oX3oVE/cn8N9v2Nxs5jLulHPlIYaRtPfmhWwh+tT1DY
NgWpkN3VDk/BEipkfZiMEuTVRy6oDagfNHWuniSpVsxzGzyDkbVt6ZtCPL8JheuKuNP6XXZCrb8j
SwtaVP+qlTEmHyT0GqGUUmabnttXwhaY5VTI1CYejSCdyM9o3/Mh28XVGgoZ2NljPjfMZNuRkvGN
h4272Q13sJF3p9abmqJLJiPtdIWlMYfFHaLFFFVBGosz5X2s+jdSnH16wbTDbtTY6znzPk8zywRr
G3e6l25jAzJeJ6+Mw+f9PDuq95gXI82Jkx13X8qqaEMXJNsKE75OmwHYxR1qU6F8dvvmnxCiAzju
7kc0VqM9P8Sdr1swdFfDomf0rCWLxmdlM56id2qojeXj3/UeU3XNG6BCV2Pk9PZP7+1q5sg8kOnv
e7/MiH3pjrZMFzOatYH/l2BTYGnQsRk4OrjVS4aWTX2xghy/49Zx6SR5YZR0FAtOX75OTwSrntD9
ba6LcnqujjB5C17tcowvOZ99aUNiYopwqsia2QKck4CmzPMOWELzsR/NqLCQQAj+UjCek640MHIQ
xZkLqrUMuG38OMUOLhAyuMWYaeawPIYDbDJeLRb1Y0Rde5gbHtUqq96gJQQsLClJ5pwIvx2s1w1C
VlJeRuMhAnIxdi8PqQNSfZGSDDK+yNKTlnEFpYDotedJvkIlhGNmF3vsQSR6uDeODLzI0CZnz/88
UyXZ8truigsRrYXe6beazbspa/kCxazqarBPjzli2Jz3xueJm4bRthZ28QfwHMik62lk4/LYQYoK
OPlxSfqA2T5GoMAufDhxfOl2lREIUp61zWr8Xfe/XYOKFuY8LkD1trYB+PGgghD4kiflkkgpMZxU
hRiijfsb3JMu7lUSAzgL6/1xionkXTPLPyfnzT6o19DjDTFtm/8wsGKOnuMZl/I2PqiZKLakFyZ/
XTuUciURmHtRriFILn2Ss7ge1P7PLTbIeUyAzQHjs+dJ03N9n8zilTrM+8Kg2ItM2pAIRdu15p4o
Xyb93kRhH0HgIhNoJXRHKNK00kPVEj9WkpngJoOOSgJFc7zSQla3MDn1ls5Ldpih038/QyIAXVkC
JDT4/wZtl7t/pUKBytZxicazuU/1ymWEewmbwxWb9OVku5iEdEiTNb3ZdSKOB1en/08ttVs70F/t
hI2+kWoCG5mol2dSNqfPmIBfI1xQJkLYSH7pH4ui9qxFs/Ga7ErWo0LB4XqLH0mR/ruhLbuU04/U
SNs+rWV6iqDwYZfqYyhUsaMINoZ11ySvqS/Cf7BmNTPuxYm9mhhT5Q+YgrjALfSuG306h656jnmy
HpuHSlRJbhCX39mU/dOLneqpPo1fuOg/rUwN6SGSf10pEuABu3RGHJzRy6fMRpKOVdKFOy4Fn34Z
cMQJLFR4oKjIoRrc3qc+1Zl8G7v+D5SwA8+M64SVyclZTX/LfTipaCWLnFh5Mb7npCYst2K4NlsZ
8T8madtC2eM94mfBtZXLlDPZfYS0QxNH1B9LWcQb+vwLxA6+fcPCLr029udnf0pxgpWMLESEFt92
CU4Uus5iTqXHxK+6TztcL+SLzSJLZBbPzycijOfgbbJcIDcz+Y/5p6QzGY21SFYDb1rrEHGMvBo2
Fuhn6xifZkOrkeiZqC+sTiRUV8bJXZAbJZsPMMgDmt+lvSss6p9xxzr32+3L0m0jIquHRgdLJkl7
qKo+XYiz0P0NNwTWL3VD5EaAnaz8FQ4X8Zesu2yVtgPx1SGu2kZanRlGK0J0AxflD2JjzyZc6ckF
HWZ/XM/GSr02raAYOe6U1HMQvikYDpu8PlFEZutbzhOfiktVT2oZX5XX+VGvuSzkupUmL824YH3e
UVjU5Ss+U5lvkl9LOaJET99Z1mZu4Xvy37uRV3EqwLGxwz+i5TDUaGF9BtIihWsYf2l9hc40rn6l
i98vHYyl070kunxuLBL8fw/c37MYZ98KlzDyqsBd+STm6NYHdZNS711XscxvYIyUKot+C2/4PCM5
R2phuej5pr0QIvuODhvkI56Iwkhs2bGiDMJw878SoyJZa53ztZxZgFO9jCWh6G+S09pwdNYRafYm
EwZ/1vxsJcREiNatACRIHkiQbokG+pzCAf4TJk9HSGtqlaI39Ftv38eGAQitOgyrRXah6MDRxC5A
VrvU9lAwFTKXvkrT/8DO4dFATuZGNh6237ifPkZsghz37H3UtErsYig485k9wOIVx0JGabIMxcLN
zjrrMTxRsrzKiVkRCaTqogE+0gksStUdzVvBJVClfKUJj2Dc4R/5pfdq4VHb4gjDcDLdbPCSTEaA
rYiLTjWP6YxM7GZiQSx0X/Kuf5shlc/nLDnskZhjG/5RP1lcWjoqpA5/R9H2mpxgBF3Qv5N0Wgd0
IrB59UemPQAJ1vDEHBTkpmwoaLWiqqfmLq1nDhv2FQ9MgMALYFnfyY43bCCuVk7nNXiWKGbnoj3F
K3gdhP1gBjLOuiph7jSuIl9vWn3L416yGIfxZj6NDeJDHeGzUtQxCkh0+NQuXHO38awqO6h5asx2
KSMRWjscrpWBjQ8eKOgHgaDZLf/3jFC2Xw1toGtICpmfCxpf+E/vLCM6mOLGNh8aXA52ytq8zMyx
CLywjeyjV7N36OdnyIYEHNNURIWTCCuw7rK5qx+Sgo190nZUXwcTPzLsrUdt+sqhVHlcK+hqi6dp
em2kH6Ngomk9Mu64cwtsFAw1qgA7kzgoIeMp4wmjondCVHRBj/A7BiklhGoJ3ABjlvav2Td999eu
gSlW0BMUI3sDYI7o/rPxu3TTa3WUhbT9XFmOqd9yYd25SCDveCSQOV623dmoXwMPMx70Rcywbfu1
eHtO/LMjQLrvVFEB1qozHiUW7lAkNF1CtjOt2J2wya4vhP5hJy5Ve76BOByJImplOA9Fl16cl/mh
A09XoG0PFPncL4eoby2TeswjfQnKINTXGE3Ev/a6JFVFILwOrNnflnGiwtOZGVfJqd9cLrOxexEJ
1SirN+HFd3XbaofoVZdtI9B5/4sloHtw1glhJAGR+c7AN0XIdBKMdJ4JUKUcvuVbZJHnWSRd9xK6
AuBi4JSSy43+Tspgi6HxwauvYOnQdJakSnX6pTNYUanTdluInMr2x/rwdWIvC7bHnouZ4NLWRwDW
yur8o84Gv/YOfLUSDgwIq5COITmtfS3fJ7jp/6CZnCatmCfKpufb8gNZrMX0xU5CtDqo+wrHs1hu
4mARzzwZoRHbMfo7cRBmY4p2Gl29BY60LpkvWdnMqvVOZXpstv+wFZOATUKIB8HYdv0Ca/Xvs9Yb
+yg9lGay9ZdbNjM94nJO//g+VZkaLP25WDwoC5J78elpUjAysDJ/z4ika2/bwp7Gax28ODpzxi4H
Uu1VqWL34JUCC/OjutUGLfQ22NROCxWYQLcy0R20uqe/YNDQD08xBz8F5lAa+oUFc/zT4X3ZGqvA
7hinbMSl5qqAawIqVbpkCvOXR9Z3QFggF5GdUwtnbj3f4LR2HD7RTVyEMQNiQqtg2ttl86BwpY0C
MHrjSW52zKSq9wVfRx/X1w7J0Yn9Nt/4u2wKvr7IGbXW3Y8RqB62enkc+OUGAsbWJ02DEuWAEMe8
wHuuT4I3eEMHxtVwUomUqJh6YmAdLDQ/UQqIhnKjT7tWB70qygogOhkVkj0bt+lJyb1xY7KZfu8l
3H1QJm/GPCUHyzgBc3rD1nmZm1Kl2TFh9KZfb6Iu3oagEiNzTmKoJrNG4oSkXoeGVPDzMK3AmfXG
Kd3v9zqWL2n02BGGEneyTl5dPYBFabpsQpOYHRnkjyho0h2Dy2mB1NLJIEbbqpYW0ek7hujDE8+B
dwrc9obE32+FJD/OWpcsViV7+Qk1D5ePrLg009ZMIhpvsKCTtR9Cs1s3fjCb5+2RS8WOCXkZOXdc
tMl+32juLbcMudft5bQ6jaDxCLLOCBy/woeXerLSz+ELIZHGKnR1vuyXyy/0x35ABauzkpjZvhZG
TYvBUl87szRLQRb26n11aT+q6c1j9vuGewwkdWa7KXz1blCEIEaDuVJAt4SKeH+pMlBrr4WIYphq
6mYLJR5OE2NjO+ehV4gqEy+VJuYCDrOg4hGvU+UEZ+w9gYzMCotAdPxjwWstjSuEUTKzpP2Sq7Hl
ddoMY/b2vE2qJ6eq+EG7LaEpzIIW0w0ILY1a+Di4//QsX7bAKODUdSMu4osGfpB4+ay+V/bqTkJr
SqMM+zhEoMDJjQqeLTtosAivPqJ8bzB5xfTpOR7vhQW9syzT0n1avhL9ug2/vojWcQ3vgCW1+1zO
TpntcmXMYWdx2wgKh/VnXGL/+IDIAUCo6X7xhV9LTXgCDhOZan0uqtYnx+hl1F2pTmqr6zh9vSWw
h6GJhOLTQM5UAc4QK6/dv7DcU9tMsU8Zju2Zu4uWD+OQPCd2NzshOb4urUMUGZbvOjNRdYzN3Fjr
OFdXDPQ5X4408E9dvjxzFMPOVo0CTLUE3mN1FM/IkP4QLUaV8Io5y5N/8K9FOIdbq8InCcNGxGaP
io0ur5zweKR16ERux6FgTZ0PAgS7fEcSw6gPFMwCNzL2ekbPdNONTQJ4CRAj5HO4faaa9HRlSy9F
6q+G2FhuTYYny23Boa6mOZKi7Qg7f9ve3jBm0i1bh5e373he9qB/JrcEaLEmHKcmhtUFaKK0RW0W
+PgVjl9qBkvNpCg2AgpEzj2IZ9MSG31NAPJGGW45JDIlwHmTz1oLdR/jbEU4ypakO6cKmJCLks2d
BfvD5F3nL2s9t41xk4dlCGI12XX7C8uvU2z5pT35YgMKPIsW0/qVQ1i4o4HfweGCoHXleRt0htCk
dwi4ESI7jg5HcOIusNLeOIw8XpWQCmBGUR7Hfh8mHE6hrCBqkpmT+N1YLKV8BInsKfr1tDzHy453
ZBFKIFckBxHrP1ubyCEQ2LbWBYKHOhugqPq/tY+Fh8oo1BB/8uGN5Ej63P/+7WNWLiY1l0/JrJtt
vV4FPIg4X5u5uQkpIRBk5Q64q4XoAazjezR+oAuaKNkhql+Ho3SexjnXxDnatVi6upnaNzz5ataf
u1BtE8JPXsryCL0rjI0eNB3LPmDr9TFdOyBCB+nSBDxEQBJWpLWUIrqqQ3K0s8YSptxfYjntMzdI
a9Yog5JCJ0Zqh5Mx0KYPR6Nssv+sdFi3UQUP+xTFNzd629FYhhcxTN6+4kkMnD9iS4MQ3j0GHxRc
iRm1pG73u5YxFFkNa1fMFj3w21Wtk0T85Qdo8G6NwlkNpne79bY7eJqkira8skbPzTXjG3nR13u2
5JpHheTSJG+yCbOdHpV3d2+MnPddAsH19uHjT/BbySVUfMgUc6pfg4/GCQ9PmpXAjm7sQJXz8goL
9SasIS/JbuHBRNC9109837tecleHIGanJn35fM+eV4+iLvDjpNUE1lVG87k1Cx4qEcsZeQ9JyJ24
5ecGCk2XTD69bMMA1Rym5Ucr1zxtqhdElqPD9rEIRj+fRvjlsIhdR10IAQ3U2lHUCRpL1R6Kmu6P
rCPMHUtt80vBq8XKV7dfMtb+nxgyc2wh1EyM7QGaoR7na04dz9NMahSE3Svn5TWjm2FzkMQDo4Jm
zXQvTh2V8EbNaT/Q3rCbJYVUOgQRxsSdXx8QBjV+zrGG4VmOAJig5GMvwtq/4qKZlQfhXDlZiFps
Mt5+rjp9GZC2ABpHiB2b7GDx2DPX7yFtqZSvpSzXoAnWtlkOikcxUZG+iDewJ3j8yh76oA54Q4l5
t3HSmJbd3ldafPCFDe8UuaMqXYNZM8JsGbIoOmDUhXGUlLuC0tO7qrf4OQ8XYOr/nUywMLaY1qPT
cGHxG1IFR/cw4lp0wdI5wTO2t6ERfbtVqEqFQ9FCbVvMQprAyYuXrzjgP21x+aBqf0xF5v2tsZzR
Dx/FrxuD8DKlZeG/qTLcpK0M2IqVH87YvpeaztfRKIby6oRc7C0KwrHSuNEiwj1w/z+GiKnakfDt
42S+Pah91yMpHM+QVCtSfDfDeXqn4FDLavyiNugQR/pdIqnadSe1ZIGTSrmKtnkZrQ1ccV3o+5Sk
57v2fUWdmNN1Bw3+yafe65uLbUZhh1agYq3KKmFzL8QZkepLXI/eOlYfTUVjzFJfvgcJpI5JRXiJ
0ZMHTBGQk0cnrQJ3yUmfB/JYN801rXPMfdow2qYMzUgiQooxif5utXDEAe4Ee5gwZx/mmBEFx1ez
8afuLItxLmwON7rg+OHBBbDGAEa57PihwDaQM2Boxr/MwoRgAnZLltBIgNyCN7DvHk5JNYQS+6n5
EAeklWCMCf/Jh+5NKY5MyDFSkP1MByCnZHU3Bez24cbASAM6yNfknziwQzOqdsQbB4xSM02PyLQs
eTiDL++jspisilutbFKwvPczMfscWXJxbk1XVxOKqr1uaMTt1mOU4xA1b4184xEPLP27c9Oh7Wwr
QUtqajkUL4tI6wyHKVGZlIs/YMJyOf4kH+cHZkeOO3Eqnr/7FCnPnVuydQm4wEwyN9aMwMqON3Aq
zLajnxSX/ltCHJFhP3qr8sfySVCnbqCsfMRnjYRDynqOV4AKU+726GhEPkJAE7l5JCrDS7+WFhee
oYcxgUaCjS8B6XzWHD6IZKgKrYHSpm+ji3CccJUqQ40kvq6JWtqJEvwx4O4wFqW6LFVnYkWsDbeA
HKVp/MXvjW4DAWCBnj9dtIbCmTIUnuRJC6dCmIi3r0s+liLwmwS0arkpwWlpcMEPFIFDQtPwQiM1
YeR/RpRI53e0W6Qwo/UFMkYA1wD/wQ8uRWUaGpcWdrAbNVKJPfF+LcKjl5YiAJPG52hzLwt3Jqhm
OH20UR7+yn49khjla6LzW8FXECx7bJq7ixhM+vhAz9Jju8A8M/TFY2HUCWPaJDuon9ATR/LjgG+6
1hE+GG73CvqBxewM0SDPsDCEL4pjc3AHDMKsx+CB0GiiUuYnw1Yb+t4Zb15mc7Qebs4gj6d2TesM
Ka/8n2/twVrcyCFePeLNiwFwjKY6DpbyvQ2XwCiKAQ2Bh0bID+TcGS8bXsVUsufYSbMNRjQ6YEPz
TPsf9vcTQGO0vtS1UCj0fJhmQ+pia6V+KAVSteN4pAym38U17wIO+FyVV96Cg3kn+5dip/q1l5Ty
l4M/N3GIa1zC+RSS32OLvVGcTXV2ctUtfqZxnHSphV718UpUTBh1pYrBns7HVaSGwyx0cED7QNot
N3+xVLNQ+uT7xZ3FJJphAVapKsGrXTTCGObqyILNpRjNtVIepPd41stHdJ74rXArczfvTdEfM8Xo
8vclIsZzxZ3ACqJDVZ2Jm917GzeZQ1l+HuyBP+MepHD78SQ1kunYw9OQk51NNX+ZBuvHJ0ewUVXx
+uFR2aavDrr1ituTAuNznR4GWm4M5kvL31dn9UmqSkYXo5DUdEpKMp1uAZefbtKeUItpfM6gAD6G
Yx/iR2qxdR3pXbfNTnjsspeqW7fxtut3XK6KLcmcxGj/KVY3HdbEkab/MvrM9+F8KJvfQ6vxPu8L
oT8/rcj2sf7NEimWf338fcUsPNVUr9K3Q8huitvatfv8IwuC8cqExS7jp0MNWJVoUQJFBCpF1xGu
71PkboOoQIqcXmvDRKGwiRkZ31lWgrDIMk3/iKDz3SD5xIc8NujqKNrfHdtaLBdowrOSrjGswlZu
PbUPXM9LHWSuwdmMydhZt4Xv3uOgZJXK1IClZ8inEuzOH549Xl1tEAH4K6qIw4X1cjEf/720nYhR
ig4Q8x4Tv1hBFXqhY96fl9ISpDsCYg1ffoejAX/cSLo2GEEyMo+B8x+kY6bhOl05UQl/CcYQz4DF
vgvR2KyBOSdsdHUv7fk8qROc1We5Z4Q6RsdQEFL3fbChAPezAWEp1bLLWPaieUmXxDdz07t6ccG4
oChz5kzd3FSUTcpUG8xEeWIapsBJm7EayWg78n2o3VaEFdaCcb+wHVmKaYOKuXHWNqOJKsx1fgp/
jwK4exRJRrgZrsvWbZs7D83nh3MxCi+9rJDZM31Z3hnTEYtluL1wusuEAugmKyhR+nZf32XDNeXa
xej181z1zrylAzJ5DpoiQ2adRGoLa7zZg2v5OgLHysstPO/lJhxpbQharOS0DjI95vdYaNbaj69J
BeyyHr7tSJ0xFKjG86PTrySakwCLdDYx7enhnallUVwWRfjqAquwfe1r+/cGhTyq39gB3m0jQRCp
vjj/Xr64X3EtxKVw46cZuhNThirbeo2wg2yx5RZ8VUJ3+o6v9Lq2Ky1Qzf9ifCql3MSLm5f8CfxI
M3SLwxz1UEL/eFUGm+bDZDUh4j2maBmz6LnON01c8fJo8gHA5NkX9nt1QHrYMCI5s01sV2BMHq4z
uZ9Kp5gcpR6yfbpdF+XBogsKzfBg3qJAgdr5ecoBdO86eXgwofZbi3q0I2vHUFxz/CZNhsdWii4p
IChCNAHL+LRkrruSEY4BLVgQ1zirRudvuyJboIXswV7JYnUqwP3BdQWJh51FqLBwGXX48jtg+Meb
xGMxUjQA1w+WQX2kpGISBVSjp4TqnAorFpATeQwlGvugdFgfZCp4qt+Ne5MJgzyq23cOUmGgs+wg
J8ZNnnes7gmR0V8kXGbaB/A49Xn/Lg466ZYAvb1JPvwwPsp30op97K4ve7+YznZnps4HnR5AN/ei
EIvJ4nVabX8YrCkhUJ9FmVRB+MQh5VkPB8mI2HRJPKT0sIMylfYe1iihrr5rGVMx4lvhENNAHLTv
7KC/21iZD5xeGWaP0yjv8irS5Z9+sslcBX/OSGkz5HDa4Yq7vZDdJ04eYKyonjqXRHAjOvLbonJZ
TDOnuI2Oii/Mw2s/3KwbEv3LARwdob5KFIpL03ljRyuMG9AugG1Vl2mdFs8yOA4eYUk1X//O0nKk
NySJGQKlSoebOlojcdbMoKhFBL6UyvHdAE+X9yuwe3qkiNJNI4D35ILfPmo6CrOy+EGZ0lGXsON/
pdlHO8TZ4hppXmOrIHbKtOmVQeAAM1FaGvfqx1vMGCXjl6Iwbrh6HGh/w7Uex4Z8XKvp7eAcDzXP
jTWhJl1ydt06d4oPH6Ovgt5ptR0CTuZKw8wwh+IZLayAZ6JigfCh5h1muh3bXwo9er0xhGegL6Zb
SWnpGlIi6cls6HvBjFPVrF+5eMQcgknLN23OiYZtZMHONc9j3XUPxclI4xgnVkxX48S32qCyw8d4
nIX+K/lKvPwLuH2phgzQtiJTMQXgyPrWcMD4Y9Wo+9z03vOQ5JpdjudWApfzUnyLnEu+fXeVpJ4C
mNu5Li0/8Hg3vFhPo8BC0OEdJb5gz31c1eqwQHJkkyOI2/GA8FrYaHIB8naQsJWsgT77bpXC7i/M
NubwA4zEnJP7IXrgSiUxbYWqxHVroE0M08CAgolt3V5EbvWgM6AEmkeKcQSmaH6mgKlQnC6U4uEb
78e5g8F6EevVgjrHKLyXJfG+034dYTBDdtO0lY3GqxXyO4Ke+aE3l4OU5hn9xmQGRMYOGrsv4Znv
FvlX3k5p/4rGj18+UtVJzt06UtUykgsWUdc2+/T4EuoHMaofS/DQ3sS0cGX79mhumQ1gmu598xre
hlDry3365+RFxQb/GtizG6lKOrvBnohGDSWHVPrBbO10huyzDij2ySbuKexdhKniyGFh6ImSu4Gf
1ONbPuE1FFnRyLhm4e9gLhwA9aiPshJlZkwmS7a2ggdYOcMDtuRreEVcQbjuTYHk/R8g75uHfyl4
xqYtYhX39PN8t1yATSoqhpqsv38jI1xh98lcpf9rJLECN1B6+DlN342P5Ev7MxDYsQz4EgBD0mYd
hmbnSCrkTkg5yc00pK5/Bam1aLubDOPSfucdbs3BmowiqEmUGrCWB8U6lU+2QP+yTLVx86VniZy0
rtT4d2edd2YPtqbhSv7O9nhqlEYddOoCqFIkclL2DHYC6m1NlAibZRrHPgPAAd5NHQdVEYrIhETJ
kvfBQRQgNUCmneS6NdfSjFyQePOIs7Cs8mhguGN6/BJYOyAr5a4JOBkYSQLbZ+ar95Zjkj9fvTwV
74NSHe4UFR5sdUXslmhi0teX48f7RS4a6D70BhLdodMNL9zdIV+8Fid6wYI/ekhMQ5F2KBerWLBE
qhBKoon/pf3ppRtc/Wyt2Gd7htKPRZVXohZUpzWlxCC57iGSTGUkvtwHd4/gPYFcXolNS32RkqlQ
l802fwYzZ9NZdrVNsjhd+K+QkMTl3omnkDFDSzogSpZOdR1Lq85N6eNa2HMjyw8Ev8DTcymNeN8o
bsKAKOLP2zznfkEtcFl0H/X6sXr19QRrsLZvaH/VYgJJMrukKZzTTeROb3YHGaUvQExb4a09JnNc
ddRduoHpa+4yyDYF548dtaZexkyyUQ/THc5hBeaC0dce58hOMJ5J4YQlijATD1aaR/RAJluozgrh
U8T86QxJXQi7XyrCoaYmVVODpEB1S5vRR0m31ynZ5TcxZObJCvGCd+7sAq+mQD4T0+xAfgbntZbP
MwxASv1uapI5R0glLrJwDnKMRD07AyoUbPv9q+YMJwHbL1qUOJj9xI4hMZnmA2h4RwrwQEW0GyjE
SnahYvdvfthfeVbr2hLwie0bUJmdgWIOrJYXSw4J3WJzxBhUzc6hQ+pA8vI4ck3XZzjiX/HT596j
U8UNGdv4KtUK33sSAlMhby8Fcewjr/lfuUdDMgTEHH1GnrFQn27ozK6xEBgZ6RZGRg+emDE1tFtx
uQfvib4jfsvOde4agd6jV/SupEBxbbMSHXsNynX18ewDg/BDHbOSJBnWZ67dlpuzCNklnag5zJAI
qNLV7YOnB9D6cyGI3jaZTzpo0diUFFrNY1J9iznXj4tbS/CiPrP0aQXIblQCobkthKamGbJFf1FP
iUXpY3bvdLMTJWOwixjXQ0A6Gd6fZuSZZRXi11Qo3eQiIytF8srG3zf/maQpUDSOYxP+nU+qJqwV
8IRu2/Nf1YZ8qgkswXgPlTTjt4tLGinSPB6h5yIjmSGLXNAj2ZVkWBOYmhEVjJVGhaOYuhWD4eFY
28bnQtRFL2dzPML0X/yjfkNQB4lOCywwg9yAaDUIrQ2odRyFcJ4aExxj/u5ngxBMnbwCPMb585pj
u/22T3dBwGSBJPHgdMzWXg7XXkrhZqKVjAHWis02vFKePczOAZHbJRJZ59y9caOJ2rw55NyvRsqm
aeUUESLR9465xg7Z/YFGCutXe0DtEo2/MG+2Leoki0tIKu7RNbUB9H0ilGQDD2gTj87jpnyOgxEY
HZ8RP77ILHOBQXr7jmONUmpsjei+7887g1sZC81Cl3YqQ3VSAqsJJKaKwaqYAibaXsSVE7f9+EHE
WPouIQo4t04Z8jN3MB1idsf2A93Z5ruFXojPi0Kko2rLt7jobzgWEcw4EAl4R63hV3IIukebLfE3
lGV9GhP7zzbqgDy/6hXdYq1NpRAp2uUpn1OrcuQtbIBmjW56dV2CermqdOnUvpMy+2tt5c57dFdu
yb+ZNRwqEzjQjsByFFFYQt4p3FuuWTlvy2OkR12jEBD7JIhJLS2tqJXajJ23uZjotegKaoMMi6xK
AwllHXNUpxKNSmc19gF6BycJaIEsVvB6bUdSR2PBT1fUljckSPl65QskFFSnmx8LJnr8Sgzdc6GA
Yev2FGJZz1z0FcepGzEntVjYILKndwfRETU6QrKjDh//X+j/5bdQRBsK2K+TfsjFUBnq/cYwH861
EfhHMlaj+eRVn078h6L73TJkiVYAUIpeFPUABjdsd6cpVn+pEYFGXQdk8+J4NvM3G4pgS3wbIgZn
dvwop+gO44L4sen/KFDuvNknzNKtOLQb46//YMR0IE5PxZcl3JdvXjLhM8Ln6UK3Hx9adkoZHJag
JOPlSBXA3lRwYQIzS+Vq9W59R0qI7F3prKnP0B7xLlvFmD8vbToZuEB88hRtbSMUGRXnmcIgUaXU
jLWA9BwVAz208vG2LQSllz5mB2057v/VRnv1UnOjBI5aG10N5R8SqGNTg8BQI+7kiwi29G2lfkYI
tODrypO0GLeYyrEB0hIcisw+fFH9luGouUlW7GJTGJ+hSn9ZTuNXr7xVAbRPZep8wIC275P84VCU
KjciLTySJpOL8vaLC//iCGSnRei1NK2h8TuDvyMhKzxYq3FIQkHxSxfBpv1OktYbPJThPhiNYQG3
TlqJzv8iToQTr020t9CMeqq5zMw/PET+Twolp8gBlFgCXu4aa+Btq0pwpPQo7O+jxt7c6A++iLKK
8zGyQvVFNWepBMhLuermU7Hk/1vaa5oBv8EcSVfrXaVAE8A417CJTtasPaWT9JX2xZIFYyqq9T6K
UeV/D10UqeAHJA/xQ+eKLOIzQ/+TmpFWAAqIF9MogtsCydpnE5uveUPzNb7aW+xqws2Aap0U8NeX
X4C9JC0pWdwpbLjvlECLfxzE0NeWN5xlj/FfJEdChyEo3WN9LjNF7s6CcAUSZBd3gAhBWJiA9Sxh
hhn8OSjBNmEtrp5hPWBDziXqJsh/mtMUdRWppySJTNQmYws8J5M/Xadru14pyYTwU1J1vfUPvs7u
Rd71Y7cdNQ5tY8OL1A1oAMGDS3SB887rk8Lyc2rFt5Ahsmf3dtGq+AzAYggzH7u269nmhGlnYWA3
ggLMwjpK/BPMgDsIV3xAKUPWkQwHK6ettXo3+5OHTe4K5Xmw61Lg4OlbkA2NYPohse5MrwNVejEW
sRJKjxhosBzOMUdjflUoWcYrmAnjb9QTLOKH663C8xf5l5Ecbb0P2tm7VaJiHkAi05YDGNxvK5/Q
zhmpD5VsTM6MIVLvjHSVghOyOPqUKhAwmPv4u5nhbjnOAV7cznuXLLjE5WR2iRcCuPqCJNNMX4Yp
mdj2ZecXpaGVMCHYO6Y0GdaMgKXntj7vX9tdf8ArZrBYjDX0kQaWg1t0DFG8pc0aqboahmYhiT7Z
K/tU+XmRV1C3M7mZmAfY7IuNHJa6q9LHjV9E86gRfrj3Gli+JohR2VqmnoN52ph7XfJTb1pUgoxe
t33hO7rGs1Xx/IbZOD43JDyUoUM3/Y6QMqO44A2pKaOw+euzhdfHIVIqwV8Ps724t0JfjcQzws6D
W57ShrTr/+D/8i+DuPM+IR7OzxJjs8y3A+kB1sXWCFV5H36UJmXhbiflz1S30vePMjMjrqpIM3sP
sIr0C7EA5jtgraAhUdaoJFnCjwrIFPBx1EFh9GIvomaDT8MMOovHqqAdBlsWp5GqpPyK37zHDT+x
rHDlSvgd2ZEsMfyEhxmRar05P4VlOodBq8alDVpLbSdGBC8vhdn+vjTXR5biag7IpS1rIvVIF32a
4VSgLib9frEOR53fPz3Pq+8tCPXWtCkVyeEB2WcnYR2HfJk4bVsTmUZ7Pl41EWYicHWLLGaksC4H
rdO9whDmGm5Dmz/Ia6tvxXFh6Xt0SeAzdxNHFnrht947W2p1oZ/RrpbNuuFebx0tVeDbPmBVqn09
K+WGe5PaYQ1xNaGwmOzVnU1W5ueRzBrwdwSKlhCxxuVJF3+4X3/28+0kMZZgVR3Xsuh1r93jnPZA
28fYmwt16/5hHP9KC8pNKJ2DPlXdJSRbuHVy1ZZ13d7YE4nA0SUDYi67Gp+iMRGN7N/QUuBp+OAB
YrJMn1McmSbc8eio3g7x8ax6oTo/dE7jh7WbQpgpGJsQA6vwWxVVmS+uRtdLrKRCCl53mbk5iiEK
yakIMpVmx9FL+PpZnRSodnjktqTKeZx2fJaToK+XKaD3UtYJXoeLIm2dC9YeyxsJIDiwhJv6DH14
wb2Jf4ZaF17E7GLFIlczvYzMUIx8bOpV5cdr+cVMWe0/v4rdT3eDRFv+6EyBFpFKaYFTfhHfEKcd
TKErF5P4RvGudUJuZwwmKRbMuC0JtQQh/0MW/gi5DLkz6y1Ei7Yi3I3yzvdCX7eJPcyyon/IefDP
dkbJ1eiysl0mfe9iGsEd3dBuXtjcKZ4n6S8AeWRT8aihLM7pnhOFatDUKXjEQNYfVvqUc70mIQbX
d42JDeUb1FCtDUCO906+NBc86Em4HlgPHHJ8UmFSFlQ7PXQmQpzTkC9eoFs0areWA9UE5HViaJ0y
Kd1PhJoFzc1aeIbFFFtrkD/Lna7nIvp42SGl+b9MyfA/X7+WbC3lOidBfT2Pnsep6jQ3EuT9kfyQ
MfM0BwqA3DxbFzig6LshE2xEQ1EDrW+3h8aGmFm2h7+p3uKw/jgjD64y9NqfCY543xpEcqAfiJKn
2MdXQFGvtD1V9ZovBuk0+mVR3R8c7PmoyqW8SJfKz0Bef8YWeIvLGuwtjsS0VxGTX0tu1LQf+gQ2
Lh85XSEsAbaE2tG3fCWjMKkAy5D1r3IOHS+6lUeB5DzfHU0QYXCRMEXs7WtHvcubOnEltjazU3Oc
yu/XzaQfZa2/lWxotgS9jiafWUtx9MWgyPg073MwoYFglMBI2hI4WTO0QfHPkt06+sxb5/4BqrcY
tp9UxqL5Sy7s774u24IXD66ZhlH5U7kEOIXSGI46I/6WlgiqrJ3GTZo0YGHiU69rYDYb26qiT5GG
e5GC7ZTBeYMNxmgUJqhkJblueSgnA2Wy/YaZOxsgi9WwCDlOQxf8zlPkTJMP0Q/NuvTFoojgGFA8
x4Idd96hQdP1pOBt47xo85O+1Nee4rpQB/8SEZSSpRYjVGWQEceixu7ZmBy5x+baExzO+4lKvAiX
iqYGqhhPflV2wzFMmFDAtH35z8VMCo7tzTJbacCt+cjpIm7g9oxjEUQ+kZIL9B05jCx4q8xTPC+T
1KOf04PTJKAZgT1Od6Vy/zaQRoacCWWxOJiSm6M3y/3yHokYtHICwRfiICwVqO3kj/8msFodwnlF
bjejzYu6+0RcfcnQTuIInjoaL/mMWuZsEqe6ipIkQzps54QZUFb5fhztZcD1yZkdXQGuJ88kHOjl
x/U+ZxB9clxX3tDlzwVvdMAkjPOxfGAn8754q6w8U+Qv2fO1xiUy0LlipYbGBmouaLywBN8O5m1o
riO3iWcsCGEfnkMoqiNSYrExYA03hgU6WgC9QANPxeo59OmTM7Fx3y13JrR3Kqb8xmMT2r26Z5p7
9zlF0AxDFR1lRSDFQBQfRvkGUNqVpMkG5w3lq4zc8m1qZfve05oVxewyAhjeq4rDe7R8ertboIGi
PM/RgduM/M2Vm7OH8E4wisab+G6CZeBmL0eP8TTaMb2ckRhgBnSvZVDpHyCgwfkKY/XBzsy2MtQK
0++tXdH/t8s6wtYPDYYJf31+dcvN4odsX3ZxYXYFpn2nELyo94CxXArbYDXluKpYGCMow0T8pXRe
YszFEQxrN8DFkoDPx1sm2qFVdz/mAv2yEpzouc96l1Nhz8VfZ56DJFANK8wDyd7lJEZS/nlNGwt+
TD6InFuQdHDcG8RBksPEqbbZx5ji4SElu+/y938sxEagDClm7Xh6E9uVx9QDmffYbZQTt/Pcv+0v
2MJRBlOcgMyYIPW9QJERHS16pFqJSou9jaUohTYZdWvi+AdUT70Yw+aXQg0w1SholO8mU+hVlY96
XU99I91/1QzvSImMBEmTki9o53pflC+l9A9HDUXjP/+ghT2xCOrlBdmZ62WusKgLqyXn+K0xOYjA
r1aeTlzkPEC0vg1lfypA41xhPMJEqpd0BrAAnhExPXCGqahoG4WzSosZ0kY4z3zQvB0XIVYyzzze
Ongxh6KiIqs7sBLeOV2DTFwWWj6+l9QJHU4GlfU+O7V5UkJRAuN4WI5ouvUSM1S9JYuxJSElt84R
JCDAgPYMqMEJ/nqseYrV5MopMA1oIgjscYoa38XwLn9dsFOhqKmdjCUnLTrSQUgTCX2TiKi1FdjL
jNWFKqyrXtrrTNlOLfN8ySNcpCTKwrG0yJ9WVg0eDJ8S1fY8ArzmKiNbfHCGOkyoixexdZxwxD4W
tvOBu45o9a0jOn5RDq87K7+8S0DS/Zs/6vvRs3Y3c12SekaRm+S6lq50KnscQaGXD8nB96IUqvmB
BOSNm9Ei5yttMZx0ujbjgM2uOyvM9HA/B+BCGK6U1SzpurUyHmBegyVkU5jWPiQYJKH+YOQUCHMD
GgjRGWlPtKiPQl9tZ42yio9+RDm7aUJXoaSERKUhN3ViqL18vN3iiwVb2Prg7ppiIaYWQu2Bwm/I
2vihqXmCWgegfyWXjla4Fi3FScwySW5teXfp8r6uvLG0OJkQg1TwCK9qA2J5DP+wSatVO8Zx+90C
K3UTNs9Z3V4TEdX9ZZZmewnLgVIwOdq4bq5GpZ0tgHC3Me6JDl9qPHT6knlWqfJ2rXwZa4qLLsR8
cBgzD7N6IV4pZOeLS9XKAfOGVHX2ptD544L2b0mga5p7Avfnp19UyedzV4o+PrBFiSlcAt8q901V
gOWfU2CxPAfkenV0JWxwfbK/bEk8W2cwnTLDanx6Ihb38F8TJAtFCJE03iZrJs/oxlONqnudNWc3
aan9SapDXCOwHJaEL5iBUO6Iywy+3D4odY/VMmup6R+r1IoIW7LRBMpQkXo/tGRoUfhRqbsB2GPZ
ERpxLG3cpuz4uILv6Fbxos/5LrW7SzEH/9XDumth4F4DNIDQ72ukyb4F66qQyPkfyEX/t7KOT2Jc
Bhn0sykY4YtGVngKW9SceWY0ImMiNEFlDrNLL1yNXLTV/3ARLhq1xHc4U9zsgYFFU4dcz29mwXAb
TBkIVog+ZpwaK0LnJv5eGpWyq5GipSA1g83Bq9cK80nPX/hkHU4e6NHGys36tqlJBCVD8bsDMGwR
pYyOf+O+fnNv40pnpDgwwatdE+mq6UBtQzUNlTpTrnPZK/GUVZvZW8tq5EnbRWxipdsuc7Wm2iUK
TlMRg+sqd9SjnNQrfY6jDz1Q4p4sFnnwYb28hce3lg8lGSccASE43dswgnxnv+k/rZBqYLzCXMUn
MDEy7c9bJP8FJurd18RVe2RUbHrJnEcfkXqyvfyiNi7+g/7g2gw4Y1MRgC9PyYVvPUs1U9EMZkph
MRn/qaF0NB24aw7UvZtDGC1xhJ7tctK8iFSG9DjOCiROYnUtU5Kg0IgORDQg6OfVn80XDnfv+aps
2EZ/SpD5MeYQ+haTO9vN43CSW5e91fc6an0R3PSgr2onQs/D/rSQATZPk94wGlAAfhcv87USoFA2
ODfiW+jnULe3PgibM4p5GIMr/ejltWip7UOCWP5/H/44OZBEgjYXonHGDDa2MnjtphkBVSxncyJv
3x0O+APv8Zmpn8nAAXTyic+bLIdqF+ApsmuhnQv52h/NtsE2sRFu5PuEd482Crvz4TGAlnKiuIVJ
dJU3k2d5Hh6DCVVVEYyehyyHzmxsg9fjhmL4hdrKUJzvBy4Y70RpQVImAkNo8X8Gpeo/qkwf6tTI
EXldbjhzD9vkpgC9YCN2hcON05LJtBMgktnMi5V6fm9r7go+SKeSSP4Dq+IlPLJ4MRyn/HxknYvc
A3a2thdjyZ57qGN7+tn1T65vq1yQ5sjQc/rT1EzTFuPBLJEgN4FL68YU0gbxFC5CG7BMvC1U5mL6
8ZW9bzMQmj5Ba4otaTxzY3EmO4BUmH6I59ZjCq05WLdoRQ0n7s9KUyHk5EGFvys3WJ2cZ/bZ/ZGT
OIrCYyRDIUvUqmSNaKFViEpPxXk0y1eEx5EoMb727ENYPGu2tl0eOBD+hahEyoi5mW5ZXqieYgii
gLspg3AwH3EhgqGmlu9x3XK2NIo+rdtIHDI9FF1K3LtHHZRAywRTMnAtRf5hYELUAkGZbeJYcRlP
n2jQv4zElPL0RnR2cw+pQFN2mgPK3CHY2TbKOI+z7Mn62dUIvRT+MgWRbYpBVblanqTmkMB64XPT
h/DoHXPDHBUjCkzJ1W/JgvdP9E/7Dj0RwiDC+rWhsxf5WIEBKnrPkJ6K1szd1vZNySX5jEPifXvR
X4dxV998gv/HQpG/z7ytRymM8bA/2klGZB9lntkv2BPDQgtd7/wfb7BaWwhtSZuYv4PIzTNRUXbw
6hQYfO9f0ZmPEUX70PHdIstIrQjHnjr51nsCpGCX+8Eg8LKeLnGk5AK+ZqyAKy7tMSO91XY2FImi
Jg1u+HQ7gUHp5VvbXufnHk9Wb58ndJ9AVQumdnXVN4jJjhe+qTtsSZ8+BFlCDfV5l81TSUF/wduD
N+37WyJ3PRSwj+ehezHeLMpaHg64QIyXgUzWIGbztDJBnjvuBzNlEL0A9voOSIGK12RNcYkVnrrD
xV8Y0kZp5mCGhbqOC/al+M780a3AFABvwh5DB8s1Mf6NqhI2aihu5ACiylN7xnHOzp9+37xdbLdq
Z47U+4GsAmNlEaENC4yGRR66Pws33ISNjQI4Jm+W/AClzXzRpJerEffw3xSQxA4faNd9tC4gA8NG
nZKPsReTtndsUhzo2Q2xvbaAqZLaNq1rMBna8bRFLtv88YkEVkOxYoIJIrVUOKbyo7j/dBApffNC
gDkn5JdP25Jp51wO0i+8DW6UGCrTEmnwZxKPCRlQVvD3E1BGRR6N20OIznsrQlj+cIe1rDIRytpw
1s3qK7s0o8PYvQlR1iu/BDtWgaVF7/It5DADQtQhJF/pxaQzM3RugB+oWctb4iWCISSO1My5u+Rh
k63TSVyJtzAX5T2OrVZ4fHhHK+EIpYV/4dUxzWxi+imY9wPgH+o1jjgJ/fhAjJNW1gibHp8WH7wS
2TRdOmJmUVZnwCVlC+Wxga/AiQmXcIA++A2uVbYP/RtytvoAKb7wuIsQ0muDyovJKQvS5ajqNmsX
KNirZwq2dPVedGfdY74fR8LlgqzMUlSw57td3DItLm6A3c2w7DuthKRFaO0nPJu6YSw4Z10ALqme
n3UiNMetjKs/nRPlcAliX/cGXgDVZjRpmVAavq881VHyZF5BBmIKXmPD+OJCSKjTbvyQDBR7jKqf
bkwXMUChO5xJpsBfQ4ropI0e5f0SKSE37TPFujbJRDrWJKIiNVBKSciXrYQhVv7m01zlbZk2ma9p
Vdawp+14hgiJsYNz6gRgVeGLwx7orFBX4kqdFaqSH8nvYN9Y4aFdNGhNGpDnxStfPXxZednFRdgc
sIetWbNKNpQY22bhPKaK1eML6j40LjVRe6FqUUJ9oelPWoXkm/ZTd0ATv2Q6xOFhJhDFcCPMvfn8
pJ9o9MpqPybGCE4qFotH5ANvipFaay2ZrVT2i/DILZfizyP+Syvflvr1o5DJxIYphPxxpfRpL0WS
UOX8ceLIOObAjTCKYIf9ZUwAvJsbHPxr/FtAyvZlUJ5t38mML+mOSw0YuUaC3o0qIj49iLPmRPD3
19gpGWh2WJCSzw40dN5FVQwXqHekDHdd6ZWRx3ewAu8AP+K61irSG1Hi6uORXjg5VFfHE2K1omb6
hs3Yht2qpimFtqjQTPLPdWxsEmlE8U7/+Ft1P3mBHZc7LJelM90S/Xb94hBiBruNrpNyfiWVHcwA
HmqqHQwtO62Kp9Ollc0WDjPLqIavcx0Skqfj7Pp57FVjg1plU99HrkIclk2Hnn7ObwljKoSGcjwW
RmDkxmtaW4/6h7/uZvG2s2dbZcMB4fVCOi0QV3dbLvsXKaB9jFnpYckOqXK1INP8E22zmP5FV8PL
6fAAmSV6Gz+6zf/oPboWqeXHvwDiEDD2TZGpl+Ub6auyK4H67Q9+gSssgwen+DL4SuUJIQwkcGgd
4llWBQwIvVHVoGsWyZF+bxlANaqQIBcxx/kz2mQM3X2zBChMb0DPFfKPgRQlVX73VRt/DLHMiCtL
7PsSZ0cUPyhJq5CcfALctNJUhyeDOkurBCiwSY7zLIXXH31D4O8frdU2e7g7v9hQUcqJJ1bUajM7
G2mNrsgmlVE5q2mMH108MLtJjXJI8VzKcXUug/sh1C1D/UNWJ6e2zRiUXJbh/s6NcwQzC86DayGv
dxAsj5ADuq+AOc6FRfnF+luQa1ZSbXeC8zU3LO+WSfEQ23UaOEnogRF19xoqKDdzbMBxu1DTwWjX
PkwJaQ3CeEp1MEEFdTNWVTTRAOv78RKBvPngz1Mmokp8sJhcMm+MWUCzALKw88HlQEbC9biQm3rC
zuP9LpUeW0I4PBrV01FzqTzXbCyXpUTGSYGEwArIxSIamOT82kNBuMM9FkYQuxVV6MwQ5f7E47ge
SiV2kYHZplasW0iJXOg0seHy2HRMOjtN4E3EwMYJVs+ipzwg/ZNqnqdWMDXBQsdx3OJUBj01unqs
YuzYzLlns0NdfOQ4xxv+uiEUSLx89qZlpXlzSCA+u8j1niFgH13871woh8w5FTeCV/yIlXGYb7PJ
xa/7ApA1lf1nwR4SVaXg8Xjfcm/HT5dLrUvb44msNbEnQiNst6S56yL4NUmAaHxflwhR2scgoJCE
/LhWmjvibmFt+sWOKEXbafAY/4vGhlUbB8gtJcaUyOH3vU1cAhCGL3eiJ/Hp62LUChJlQuyUvAM0
AsTSW2hMOfGoYbkLfVrZdFsGg+KkGGTMz61YBmvivXc3vhr2eviD+XUtScQ62JZJhUE9sRtsJx2V
uOP7xiZ8yRWBhlGOBnhAnSiXUN+R/I0c7TmbmfC+o6VbEJOb6l9dpaYHM2uwK7KRwurXhTdb6JE5
wvlgB0XsWIAIvKw9yJTJbasCLRlWSYJVpvrtxAlvK79zY3n+SW8F8O3BaR6OLlhR+W4Lh33kN90P
p/rsGcaAAuK3b/L4EQKg1py2XwcWuhiT6Q962rkG2NUVyueN62wbB1Vx/XdH58ttoLmr88DuLLqX
HsLQSYkSlYo+IcGJZvuttpZz5bPkwDdqobL0zzr7aYgPOO/AhRtUJC8meuX6dPxXBOYfl3oHnkRj
33GvoWkRar8Dw7jFXGAfD+GZSwAbEMJ6LwflZfcJbTC5KBCb36tPTC6Znh+JQmmWzs43DZCgCbl8
DzbV9SgKN7q3Ew8dJbk3MsxZnuWbhL447nCx0IkdWNdURx2PGC6Y3lSwUFdzMDQnTAXAUDfwSdS+
XfWHlbxGbWWE+tzwP+1NiL68s1Cz1QjrvAL+JJYCZbVPEoGSUjSTazTTlVLp2YcCcqvjRSKrEX33
lqSF87PVb+SVUm+r1VVT8RWFmiIFmXM/BBSG9Vde/OL1uE3IUV0/tZvyL1pJBNPMRhY+ohpSWWn6
Fv22IzUpy9DknmFeQkOFT1GuJ1GvNT+Nfvblf3mTJ7hdaz9XVBJureGlRHlvhqUFluTvH2tgnKqM
SkfySdfFFv01yWOJhfQ6EJgFbwg/8fm7prKzqY2+9cjtN3dqk9VJ8SPGo9CgBzOk6tMlNkhI74f6
KvN0KKPCy/Y3HbyM/LIcjTCGF9oTtDyHVtAKbTEawp5nW6iwmga0VUT+FiRl5MbI65XUWLFOlVck
IfPw5X2xomep6lEln59Wjagc88IxNv13Vobq8PoSxxvZ4u9pV8MjvSFWdNxGn+OGDkKcx3S/JcZA
OmSBehGP0l8cttRzlAb5VFOcIP63P8DjpsS93qeOc6bO1h8RdymInvXtzGxL/OPzQEdn9HL9E7zx
BEu0LiXPXdXqypslhAj0X991/OiWjx1oxLN0QYhmUpg4pV5ya4dhOREd/19UfLV/22bx/JLWp/pd
Sb6+O9KBpzintczSd6ZoKpRD7sU7nGbS0TLbtXEE5kPGG0kKLecDwjbMctu3rYENcDNAdAT+OivF
XaBd6z0oalqsstv+VBa14cyB93iVctsK9DCoz5XI9bariZ9RsJ72MDQHr9yQI8a/tmSn6vNae35L
ZJsnGoYf5/23bMfsQPV0jWmM5CActVVmvwiqOD/J/YpjaFImtZGiZ6zUNfi8yDWH3pwGdsuXP6+o
5kXnhsTAi8HE/klfSzbAPZ9c6hXHadx7UAYPibDUaAelS2dQQZ/gXBJkhl+nUUFOPVls3mL/Yoyz
z0vLDshacr2x9j06PlrwLYbPv3Z7GtWJpHQzzGlbaLzAI1Q1mAzoQjw9qtHWRnzGveqVhaH3/zPK
dxqB1Lwfm66W1i345Q4r4yQIU01WXi1LhcqYE/bIYdXd9+jIyLDiXgfPYvrbiIItakDNZgbhXAAm
8lAQSCSJ7C8pumJ8idSJhUnbJIo+/+XKUc3J4h0NUPAJ8IlH4RYfL9ukAA9TDmWur1wVMUnJtBPq
3JRcoKSPGY3q95fjIoVwEIT+HPIZ2zf+cyrQ5mP/B5nuPK5UB+tl3XUMDqHn1ciNhdd/iSYCu+AP
CzmUDgHD4ppryTMQoDiwO85qY3fp2HMIlTS3Y+s9qy0SSSP0vc/KNKrcQ/OiFfgiDxczVuQd87Zj
3OoyotGuqnqDEmP8NwRJhNLoXlDsutPcFfxm0CwSUtJRNK/V7cvGWSJSCxCR4FWYCJqeGy5PmiKL
73m2S3MfX/peReeOKin4z9vTR3d7x/JP+cPMvKnLMPzOSS4TDySf8aMTIgYDbtYPkf2zPTHV52Tn
WbF+EPZ7p5oHvsDeMJAEcx26KgB0/6oTY1tdRM3YUNa68/ybHXrrl87x7N/59lNo5ptylW25gL+l
gGDqe9q7M5IaAeRGFnno4YRiFn3mmQWhqAPO7QtOEqwt3i71QRtGuTXaM4zw9GQOipDMGUi7CQNY
zPJO/3pSRtD8bTdGUszxePst/8LmxgIq0MxKm4vSi4GOMXpovN1RcKQVEMj8aqOWvX7boTLbZ5W0
MjoiImbfG5YE89Hj3N3G0U3msel7RAgWzOhjwjCwzpRUOWfAec7qeFoeD9d1d+jIexJjPRn9IgHl
1dS/khU7YrFscpVG/xRnNotN+oh7kNkQPsqsgGJhPNvOrm06SfMRURav/78wjA4SaAwcHrtjMLt3
1hUiMCGCp2jTuNOWaxRp5g2MU0q8xS16K7+EkGyiDXyz9JGDRGiK32CoVmc0dFqnPDPjeAEelh2+
S/qvM8TSjr+gKaXJtRE0soixcWKWtirybn/AqurdeOwx0dO+vwWjrRR4HWypQ3FOTgsGZZP7RbCz
8/gbFIVAG3fWzPm/4CaqBn8Siru88hdM1jbtqS97JeqycuUMu/QkmU0r+St0y4dF2D6ChThNjHp1
CL33lHdSnSady/hJ8JlB2oVS9AnYEsuVWit/MT7WTKXMqxcSlXEZjyHq5Kx1t4Od6r1othpnEIvV
uf4N8NsbFftEnzE+yMde23j81vB4gVJfwbZh9uCbltBHE5rmainB4aMoZfF6vQGs2sgSQ8MbG0u+
xHgeXFm6VTfr64UkwYdQiBVdSQZ98QnqGLDBrvMRxPqslwXBmxxyagmPfPMpjPGgqMjZp7FhFfeB
vmLxmk9Uo93WpVvJXwE9sjxJ1GbEIlSORHNvwF7/TdY3dbAoqYAG0Rkbd6zwHm8zZjbXP/118R2J
uYpBT0sAp4NayXapTkf6elePsK8dcRvnKdXVYpgPNdwUBFiJH/T5vrmLgc8+Gh5USBlDzyXQX2k8
pxKaGTbYN9b8k77mVPq7T7507d9e80pb9LvFn/Nt9T17itkGue6FPZe+3YrWC4Jn4pMj3PWY50Z4
VdYLTh3cj1gbwItZZjyX+9NMfsb8egXSlTw/EaCVBavGid/S8pbtqvt9Gma80ClvpFP9eiXN++D3
TDosz6VV3rHiZ4BZCA0q9ic1s40kVXLqgv2EWmeR4jX7Y3Mr5asS1MpZ89t5AT6hBMFpolWFLT2o
AEHz/XHImYW7f62neqWve1YWO0ZAjfUazv5sYIxqoW9lbaHfYNbxwUg521l8oHTyaePcRXZO7ZWY
DgPrA1ZTp12r8WUASrB6tO1mZW4aGzfPl1qIdRnKU/1SyYXv6NKawqv1UNlJVWou8QC4+xfKm3nY
IYgYraIYymjLnA8Pz1upFSzImu2IxfxADpdbAwQSIXcZlDx/YZbeiRF4pfpLs1XWiRcRXQl0/BR8
cnSlQCYlsK7sDc8PWPFIJ8OHy3GVTNBVIo2VLWrjaN1M1PV9odHFgLTanmcTuadpPks/uV3kWl2j
7jOsfelmYkng/IivA0I8hwhPyubD23lKAlhcxpNfPnNMhjZ4oXiMiaICKDpjv3HZ64WWFUtwnbxs
pqEUWm23+kM5hXTAyvOn+ILqiXtR+Ey3340qrOuXgaHAy/ExdZKdlF7xTRI7XOTHeqDCNZsVTHQw
Ubr252GWBpXb+ZVTs6vKosMT1lIbDYbme1hfgjMnpNkRuhkJ72Zw8tGS6rHOW9S0bV+UO1Vp0mfA
X1a5X+vg762elktXa5Q0fdHGUZTiP8mtCA+AEDHlBJ88myRbRg8vFlNN8z9ETGWdvCZE8CRSE/GW
3DLLmohdCRWAVbhajH5Ly/VZzXRtUMhJkxd9t4l4sbIoy5utQ94OOUpi5O4GoCt2UBDEHOqI+DS3
eZEi20eEWUv9oEARvK+19zjGvr3eWxu5EpiTtoOEA0hWAbM65kaBeUYXjwa6MFhdRQ/N8N2cYbt7
Nyg622a9T5wWxlTa6b87P+IqMmYX3/jJFWS1ch6+MTUkyig7o84NNfKFl+cb57/4vp9OTla11DAn
up/MGx2oNhq7zWbRuEzDtumbx8oJ+tAbQ38k62gdmuZN2a9q3hUEAJCmSDbwLzdPF05qdWFzpH+m
fb1nv/ZG/UX3wRYkSHVSSCqxSzX3U2s83Avfs8vxhczRQ9ZZ3FRn76BLuqgOHLyVQUNxmXXDquLn
se5TEsYVx3hFCeV7V3n7YB8mepvap25/Xwox0UKGS/KVBSluJuBYjTlIImPL/kAb6Pf7dXm6wNCb
LUXLSQ96DeGytoLgy4VAhxdchkpzCL67n501p6ThrEM7z+divNOF2MmpMrKeDpBQfWh9O7LatLOG
aSjgMsDo/2K39K5QNq6jKmN1cT5vIJ5C4c/1SnX+ICkFhLPJNvUb13nOfebYS3RSAfSfF2wnnlvh
w0FXUfd6wve6K3SzA1GNhUNjOb/MjeIAQMj4EUeEoPLb5ri+qV6gHXfNtwPWXfh02anWMKlYye7j
mtNruiNTX2heMs2E04Ei0+vMGQOTsXs8O6139nK0yBm+2NfW1wKQrfgCbTq8zf4LnDqhXzpqmLpF
k+PlcXNJJXmT1OO+HoCYco64YNzMGSfrT+EIzmiTMvYBEjuKqeQJCVWpl/UJAZclJGVBbLqc+1HJ
yVg2BUO09BvoUmgCzcbkq/9F+oxQTo32NOHst100LrOtUjzubtpbjjl48HlCmSk5l5obLHdHG/ES
2sAGGZQeRQxWeEa+nejQ/SZo2NIsiSH9C7rCCeQUcGG5QtZeE9uX/9pfjEVgnaxRX3jDGN1vLsCY
A8Hzsajg6lntcW/M8d4xMu//NW2vv0ixgzChMhV/UDhhTpTB4Fpdk3sYs4+daR1cz8ogylHNnCnx
/po9R3r4+718/SGfYFLF5hpcN5iv7i2mFtwohiVQHABCTKgom4NSlnKSpM+uweh3mddBHUO1uJIB
h9slwc9mzNU4qImvuqRm9hUmpsZ2rRTR1q8auR7ykmPetFMzuBMN1OBsfQ+kWa4mncJ3gPXlKl4N
Z3ym14eYT4Ge+dRM21g4nPkovZd556dqhk77un3VkohqScszKF8C7gHRRpY/eC41Jovv78n/KaNd
mQbuDsGzbz3N08snKs5jgaV9HmTP294l2Jhn3ErhWG46sYxgjPkKlQx1efUx7ZNgD1t7qTxtNCam
5Kst85mkiRhC9pJGP5dy76JWrWtld3caKGm2qukGr1dvwIQf1JYbKIk6Nb88p3PG3CWw8Jidhsl+
8cU+mB668b8MJEORHXLu9wXhhGEGzCZY5My6D4dDtYCCIyuYdq7IC7P5ukJtZDREX8Inj76e+uJy
oHUTlIQtnyXusLpVBKyCFty14Fyi41qieGlc4/JHd2yNZ6zwW4JE8Y13fuoj//xSiBx9+s/MfLI2
3jkb2s90/lQyf9ljR5stGrKXaB/l+x0C3cnpe3oui38KXdeTpTj31mV4InCUCSF7w4nBh1HA9bAj
7nqgW5tJxQ3UpKm0VzMvG6zVNC6PimjgbU1D8RsOJgfjm1UHyxqKuNL3zRN47i1WYMZvbfFkxyeN
3h3w6BufUmT01XdCJbuXwWvtXcLSit+0tbKln+cssAytxkWG96Y02yb079u0gLUirbDkdW1twraw
MK+ldOB4itR0O0q9mtroWVvpKhlVxe0s7a8FSt8Y5hzJZBJQm9k5UJqvzJYg72VLPapy5K/n+DFC
FqNfW7zyIlPq5O7MPsPbISV2rMSgYWQ8uH7W+xPAgArKXHeB8pHl0ATYASDvqNvBRo8K19fJSdSh
3ih9y/xnCdnjP7ZQo+O0cl6J+f4DRtIknm+9qKvGRAVH6jIRkfZ9Z8A4fwBTdb6iZU3l450OwDr0
j4rPLowYjlrWOSNMtfP7W2sPjVO4tdAvDEBsfFYyfLkjvDBssFYlRiA7W/kyuKw/N+NC3sXlH9vw
vYatx9ZZlKw2CwXyaYB6JwhHdoRoZuzFuPYwRZlgjXn6Jk1naOR8rg5GWsm7oZPjS4Bb4iGZn4Ld
cbBp9PWHNz9MpEAgfMKHvAB1iZZgRt4mqW0FfEOEtVURxpMvHldMJCPU8hRh7VZRNLzBX99M4gMm
9PvDe0d9V57/HeS8zGxTKYrMQfxpWw/jtF8vDITQhqg47c2/hOgyASSKFk8RWMD8knlwtFTcRjBw
JvSnKMY2ntSLeserTOVH9Oy/lM+KKw4swj+OSwm4Uy58bqh3sNqfp4T+HI1HmFXo1Uje0Ef+1kFZ
zgmUl8c0ffGNilUAsyw/Hzi/8K/eJG7UigbyzxzG3z/0HU4p3O9PIjnABiA3AU7LNc5O4r7EQtqP
eLKVAQluPDTzfZBSB6Vi5JKTrm93ZhnSP2ag00UCxSgEew6O1NyH/Je6gQjre5y3+WRwa0YdC6bx
1za5bRD4jdOsShKjNdlIMHYO9bMqhU8uBfo14Q9XNAcSYzodzOW/Q4fNjK7XAUR+ut37lt2coPDi
mB1td/WDZRpSMbM50on33iENkxmK1ALDsxqqh57LdxacfoI/rMtWccgLmaQjAl8w3F1O4WGvaR4b
o6PvwCe0DJ/L5MDeR0C40FIEZ4u8d5ShMwz7W+X6H6sxLVhpv4Fmob8EOH2Ms5wEEs+h425y0FnU
j6apvf8zbRZlxi5FmTYpMYPAAjXN1T+mLHPG28si/La0Q+CTJwUXfO1GiTGNb4vspGHSSjP16siR
3VhrhasHMZRkXZPbC3G+76J6HhJ4oRFdAvbHSK/vaety3hAxY3VU6GxJDN6+pkL4R2GOhzWkWvhR
mv/JEZ9T/SoGsAJb1nWh1c8OG1trFcTkrMiOzsu3m6mh/6hkvWROwKH/KlLLveSV9Lx/l6lJaaMQ
uP876jrvCXdxIqUVo4aF0/g3Q3F7Ta4FFWcZ0xaela6PR3sSxacsqAm3+L4FbAvwWv6lhOl0M9+W
i8wb6qSiaCqDsQvm2pxrf0/ls9yy7fkRRSaqSAXeT/ax9cvibSc9YicsuuDkwhXB8z5HULM0zKd7
KOPDDkAcMrXVo5cNdf9NEF/Y5W6FDZWKRqdLlepmUDoa1jzg2hzRDzVMNlBkzQItGtMtKF4PqL2E
DcuUbBkXZ9TFr5kZEhzualJs9gAEVa9/mhK/3twEH3EZ3oqfM75Wg2icH3r4HaEXinuHzOPg4wJd
51cYZEjnrv320UzIg41D5B8+cmRPeczLAFxtz7KiXuXvP8lVkl4oBX0LaiAXzHDRQ+KKvXGLoxKO
k2qEsKVLRerZBEQYt1L3K24lgfXckRPiqVM3nJndifv3XpFBl4y3BlexEzYsRaRuPcJhSqmBNpDH
9W0FAbHwxTZhnu7zQfD9djHf1mH4RjMVdrkJ0ZHig8qyNihiMA3pInsgSed1/bNaPj8vXx0IsUzX
k4g5fZAXGKOE+yCVqmrhUDtoHjE5+Ir2QPDNR8TS035ksitlXw8hi9aOkrosSv9aF2bNtLmYA5bS
xb48EW2wXlP741N8Pm2vU4aT6fBXGbp5myEEMw2QD9Zw2GlW9ILUfP3jemc461vGlotr8n9Ix0eL
VDDVtV6zC8dJ1XQV7sDE2HJHOzsrzaf8ES8AufrdejGb2xGK0C65U+lXaPRO3LEKTLG8K1ZkfPJ7
JMAQ4Na4aXAW6Q3t+PNDj6H3gQCKxajUWKazkErvKeHxqWa52Zt2zan6mwfME/+3HI/yL6wqbm2y
Kix14BUMOZSqxgeMEo7cUzVh9xPRj2iZd87GYBxrC8LRiGTEbKK0YZc5nsA3O7zKxNiq1H0lK1D3
sK7ckmtMBBFyfJ6nFw1kHyHjotHMhCkAnrIFy0gVTloz9dDcsf+GdXdhbO7QrZhBuTTlEnVblzU9
TlsbaOwvCWwZAPPogL+6WiDJmRLYCkN8L0AmqBtWD6Snw6sjt+QLQ9iZYatoZf1RV7SPDaJqLT2N
//euqirsv//uqt6Pqxy2rpnbRI7X5Xi84BLrTiNyNv6VHxdyc/nZPgD77WShXoKtTx6694BpQCLw
gtbbevraFhX0ZODmq11po7V3ENzkteMyL+meD8DLB7Yl1HG9+XSAe0Q373XZKQGU+vvrOeRgheAd
Ysfyf6fKlb74rncHrG2oUhjX4w+wwBLKsdwdcuBaAWfE00CJJ3SiOCA6SEHNGnkz2Q8YoE3vi44U
aKEFmAMCDBak5oqX1GaPd1V7WNQqTP/6Uo1h2wGy0hyRTgPd9RPY/yXi7hyAhcYzd2pFW7zqJt4Z
72GPxmt3ssdWzh9IfZvu4999CMoSPLlUKSuivTgffI/5z4RFFlcFZMvvUOUlnI+Eta63LqvUxvJu
oObtx9/jXVL8tOE2SUn3xBGsGkCnBNgXOmeozTf9Mo9sSAREfhI4tfsxosvnnefJgzxA08UHoNVN
06miMsuAmMkVp5qQRIyhpCYl272VMBYb60C//XBkFMh9r+iIyqE5Kine6wqsFmy6hVJcA0U1dEC5
scozUbVK6HEJBH75hdcyIZ8uMuXvXJmJB++tl7d5Gozn4HX2djcaOkKpQrImpPgcaVTxco79vstZ
hBnaA6UgQBlWP9OI8op6106ZiSsoqgUy7lVTQTeDHCVZrJ6YPp9GMBsgvSxiHV/Rp5Md70ZTy04W
dywKRZun8egtH3+5BXWpU4ZP+9AESqJoKjknBg/a2SMoJoekqCZCn7saurFpjZnWVlEt6AMU8Gbe
uAGYj5/duh7rCNr4tMRJhMtOM8xXqQwf9J4xwKFihRUMdV7zULJlAxz729cqhZF5qcmlc/NX6+9G
Pcbx7mqnz++cEXFwxQGsJZrHY2InQDXfXB0wa5ZMQeUey0klJnS4pArFfDvKBm8qgr0jTzd/u7Hj
wyo8/hBnSe3JMAOxaqn/lmoTxJphcgMzM0LkuUgyocU3/gjedZUiUSIhqjsbxHexhi/msO675ZOU
1u43SgRIUimMTeHadhygOyX9L7gZ0Kc89Tk3z5yPY28yXY2eIpVR5vhYhaIf5tUYYbSButlu900I
d3t8sdw/3Vsr7DeWTOFhWKBt8IsOmMw91soNqVBsf6mXdQRmzs36Tu2qGwovb0p/71oo2aX2yqi3
zXdhIjIL37XmaO03WMXSKsauLoDdMN8pe3eiBuFy3iM6xNNhmL7xhRg9asgC9DhgmQEto9/g75AK
FnD+1lQ0ZLhB3NQcnXpp74oRD0WnwKQnqmOKoh2Y1VZ2j4ULZLk8ddVCpFVcF856qwcr0LlE6SKw
MW3EDbnu5lvKUJlJE6IJQrXBThZydPLIl5oMeVLacKs7huCOaIlTolNAQzVGPNTN6MyRmO5T1V8X
quEXsqAe2roO8jN4aJFZRbq1TUgO8Nbcuv7+G2oCYj8A2Tbl2lWxSUMpo6eZo6BRdioIG2iRPOhO
Ud75xQR7a0PY05iLyt2G2AzOOadBz6YzVKUZCUbzl6ZuoFKg4CJi+xQ/q0lRD9JNAvClYNmsi2en
CaFcVH2MNDs8pDqKFJEnSpXjdkI0iz1L/yRdQCLLndTdipUiOKv7+49h89ZKpN+ejTc2pHOKLSOF
AFhGMgtf1hLmUqHsrIYF5YOQdFkV/645pDnJmCizFgDpQ3u56zbgHJGxuNOl9qM14x9SO8S4cNxg
ax0VSAvec9er/egM84PxJKyX33g8eOnrwwJRHQs9RgpQVsmJYTTQHUdvC8pormTBJ7eDyw4gokCt
RWuuW1th8mgZsw5e2eiWAcDhzLwv0FRQ1TAiEykPyQLD+gqrQ398zIdJK2iq4RELLy5zuJsNtfYQ
aJjtHL4kILJ+O4KmIPuh2H61oYNGDCEbPAiSjjtfKVcwL4/hvX8cTzu5xPTzu83cOYT35XFDOcIN
L1nxZVxjmBJ7IEhL/lhO2EmpyIVyr437Xt9mFBmI9wDY0sLToXi1223PqkBhWuIW63pbIYB/NAc4
W/gq5O55YmfPQZtkfjnw7ZvF3Zza1hhCkPViF0hi1Vna9g4E9Au1KGeyue09k70o4UnEieEgloji
UD15vyhoIJL/Y+7/4otPOyLrwKuHnolRDfv0nz6050aCDAIbRaKSYigLCHxLtQOwFN4KHVFVaMvI
QKAoiROMwq8JoSJRqD/Ps/HqUjVuVOnYZpZ0N2f5OCQ+BMGaGPbYZDMGoaDEus0LoKJ/2RnqW3xT
+kB0y2yAUXyGBu0frxonQy4ACfXf6zN/UrX069plW2jy0vCie+m7OdMd33mj6v5IVB5D2uYkp2bi
gHXdJIlZ9NPn+wrttLqjTusp9rzsyzQs/mBDnvuxAhCRrGib4eDscJvmOJN/0Lj23bunI3A2XIPd
yEuORVKo9QzPDwvrHT64u/Np8847GfqEOaJpl02Q8ThrzQGuWxltqcOodtwSdKJGuh23uSHTQO6q
Z+LYS+Y/mASgbEVz9YZk1XRq6iWkKge9Yfxs66cNoNw0i3mIOo/0qGdQ5yHkF02BoNyC20KXQ38i
apg3xkQ3ObLJ7Xte3kPrT+q7UUDj4+E8fLuQ/A85mNcewr+VurppuaQDI7yJM/a/z03ZbPf06lks
jjkKlrhpYVSfyQ+R5Pg4FCid8250rZizkcKFqyKamWomOaVf/j47YPn0SlV5mnSw46LSWFIndzRw
rqBgJe4Yo1xYtCoQ/IXedOrGpyAUqGAjq6ZG9pSgu1Ri33ysDGLk65xV98kRQCKoC8CJDZAJANls
huoJ7Q/QP2sXMMAm1JSSGJ0TEHD5eqW168GwozwIH3hzyWrcx4jFMgCXiDEeIXME639xzrS3GVZX
DPMeHY13taGTRfJ9ZtnocWlgOJ1vyZxUPA0Hhvs4FpderC++z17FmVHprfLcUmu+xJhVfnre2O3C
6gpVAZfdjYXFh7+KUbEPsehOfo9dgU7iZh5YyQsLAqznXGHJaIZ5S8stwSQdacvdtWTzXzljMlfL
MlsUpTDu5WXZ03wvRUVlglHYd8ZI6cd5VHZb+Phu8vGXXakxlpzA5uy80vAJ4e+qfEbKgSGM/eAV
9uOrs9HX3zsL76S2YE2LUoGAenC5Fc9NyutprCkRE1T2CnbSyJGnYvTsDbs5K/i4cd+Zg+H8MDGW
zKEYSVUch/C6F4b8+6P1Lm0iklZrm97v3dgubAijKpplkeCYBzvDa9RpHZHEV63cDUyaSDL/M0TK
8tlYYtCf8Qk7om5D2d2JAVdo7dlNsGfI1wU6815Ts0PkP7cDwrGPHde9wxGe4oLhIoOcNvA9dzhA
kiZBN+7LFq5ZugHiIqme7LId/ZREXPM5N1QilJfGEcswPc2ieT9l0M/YNjy3aChWP/IOWRmQ6QZ8
xiZ1Z+HcGJyiVfDJI3eC9yAWLCx0ayrJpcPUOuNLs2fqWmDVjc4CU0bHjF+V5Ur70VOiO4J7Yc6H
ydhqYWreBpeTstIqrS9MPlMFvdVKLsyMqnyPWnD/S0cL55/30k04UbqgaCJOMIZj6qSH4jI8KBiC
KF/YaE4jh6NmQNOPy7Mu0ie3Y6kFzmceYTk/bCmN27LgkHobgigdDjbzCSxA0HKVv4EtRPquDmtQ
/u3QD+O61qVpMQ3gbbHZmSwDOj9fD0f9GWwEyEULD+5JGTNoAx5lKfeatr9n4+DvBbeVSB9Cmnpg
hBl0XMcU5b9ru6lLR5uYn6Mj9j1n1CznpGvjnrddsu68cbpKgagE1Zx1T1UZHLCBa4g0CXh/6rkd
VLfXzFkEdwtWHCM1+r27Xppv9YTE/C4sbrqGDWAS6/l+5noBRT6uVAWwKQuYITopDrnuc67p+6LJ
Jx/BMkqeEfpfC25nOfjQkHSRlikUO4azGVb/1cNERotTROBIHAKzBqlTTT7NnAINCve2pQOv66pA
pMXgsBGXEeEzoM9YMEX8GwTKofjKLE1Cx8+pw739vcDQ6dSmMocvqHVeyFPl9rLm/27uFpO53mHx
8JYMS0q+RVgz4uC2DtAAO1sPDpBOq5ERO48DLd6i0QIsc71O2aXxzHTGX/llrSiKUQiqd29l4tBR
ZQUpdNJCUwHvuuipMqWXG7hYP/ipmhvSrzYLQloofN9GN9LACdiIWjr/6PkS/hO3zmhagZIoocYG
xWE78Qccy+NjeT/FFOMJ0zwFH02MJD41OoIdzBiLyvs++CgbYH5LpHrt8mVw6pbvqd7YmLf7kXAX
otZpvsKJte3+OUqMYx3pnaemZ4o29RG8RK7xfT7x295g2gXwWqwVE5BeR/9P8+Bh/ctY4V7LuqAR
oHd2gsUHNNWJP8yCEhUx5chpCISE/5Ss7e+FHLynl18uxLom6T9GRfOWYqr/DwyBOBn5UaX+F/pn
KuPs+Vihlo11JIMyBvJsHwqeCQqEJpHTYRTAdQ9TsmyNPPVcuIP+VxBvuMehoWe12cmlA1yANByg
0O0aRJwkDwbCs8JVi/CNT3H2M9aNAJQgIPktdNCjOhlY/zZ1knvn9mAVfOGfDdBQ2BRCntHequ8C
pv45sBXzF3OpKz9KbItl73reUlYteWCi/7RQSOr+aYcFDFLKmVaas+PxfcHRuV82LfvmZC0bBP++
rDOQhdDPXVU1aOM+u/Wm39d7kR7mQlLDxtLJgz7HIpXeXj2byAy/L7QWaOZao53MRZZPmgcoBFPe
fVFpgha2wYz4gco77h71+vXihekpBxBRu5gsTnpHEIf1dBq1okYtsVIiFU6d8PvWd08LAfzgc8z1
2K0gQ3vN2MrLluGytfuFPeY7525C5RMVjl7k8DEgWlP8dafvqDiSRk1Anejgfv4LopsWapQ0alVG
BPVXy8l22ujua/S0dkeJUzgXWF0eVGOfxfyqsnn233gt9ZuZYBYEAWql8HeVffwrV4miJrZabX76
pLVZQdG9rs2RPkAQktalo3sJggcziBuggp5bbRP3Xz00Pwg6zN4KUM2DVq/QSKGL2F04z3xTRINU
nhwWSBk76iETSrhDTbAIZf6L23SWDLLx0ObBdHnztKsRp8IFBTvey2dVLb0rcdSgcBZ1gSgLN3AU
RefPPWjvHMhsB0nEt5bLIrp1N17LqBaE3cmxJaNg+AlpjLcYxqeko0nSiE6U8VKgSNJxXwN5kr3E
EFWuiNCAD/zUt7FhZo64hD7qmW0zObl2V+jJgiK/t7IGH45lZJ4E6yB36dMzjP5iIuasVfdnfgcz
+MZsOqs74WnHuPAg73UKtlWJq/B3hXeYngf4XiG3gm8jF1OIjRQENk3R456Op5/ZmvbJyDxKTxEu
pIOiKjffvVyfn2HACyEzS5Sn0oztvHJPs9w/JjmZpKnjAaQ5IRN2K33T6GSAkFou4gHzwx/QWYx8
LhvHPjs5Kzj+CD9+Mzj13j7MWgXjH7yeCrapoZcES7xWSqb5xOrHnkiVun6C98duf0hyqKS3vzO3
KYAbzjfYp+dW1HX3aou7VPqN/ZYqM5beRhP1eGoymPQ4BbUWii6ueYwA79zKRmCqVYsZXawGqdI3
tGukhuxFGmBLhIyWpdRJdlcxuJHKVCWzvQFTmaijmNHDYeKmUNiGiYuSxWi1S2CdhSYR3IRN3925
CrNqEqEImH7cFhzXfK2VYvxFpRAX8Z3CdM19QjJptim9J/iX3Lc0wuixBaqy1JK64cB++4gAICiq
R/buFT0M5JNSoythYkvsMhL415Esko6YLXZ2od5Ii5wzSovDTSiQwQmVFxOZtEgQ6AGDD2DB1aYN
EEIidujEbeoljODpnl4ywOe8pkVol5UnfEwgUbQIZCx9tvRV+SmObxF1WOgI4ypfkHno28lvyEFj
ue3hh7rLbUrZerCnq+TmwCyHZBk/bqvGXClHb3OyUo+VQcFD/HlWXXimRkpdovFt+2rPQqLewD+f
PSmKBAbi+sCFp5JWo0GwM7bpd04BC2xs+vX6y8//QCCrnROLDam1rBSd7+bAde/uKFN3FUiy43qf
NRQENWZgPq75UrGmo324J7egXnd3aOIrsnZDzWaFRHEvfFXadjnETqOJJTQ7ri4Yf6mVVzIVQKPo
T6xCkEswcYj0r/Coqng1erUo8hd9CEOKLPC3NMuwa48J7pE/uPHEyMUdCPGf0jKmVbOWXA1+f6wT
cDSD/HeeP0zo7NqmyCwAzEh62Wd5wa8aXQk3XChxEL+kQ3KLp5aLSHL2uPt0IyWtDiPet+ZiDU2x
jqNNVdd0CcnVx/02rubSR6s79+VwTGwL04/EB172gdceXoASsLK592haMdpwcIzQ+OVnhD2ALg6F
Hhc2UaHdtCYki3JS6Ga4BY2T1czujDYqsfWhUcUOfBAaTeikKBdW1TpAJ6F6FOqgnP4fxIQ4M1ll
xDUXizAtMlLp0wlDaT7YX2yRx9AR4MaiSorhbScdZnaOWbDgz9m6XKcvSE9XksxjWpcqk8zIxKb4
RarTs5vrX5WGVncqMNTcodSSiobeaVOtjljf+Bn2bpaWLO/Ua2+QtHgrz5u2FZamHKvmU3oQGwev
zUODqMuz14fLHbZRUmXz8CzZpUIS1OizEl0PYMCGVX/MbmRHRB3euFWlUFzRiViFohRJS2YQwAAu
+ZJIrU/FT6OtzjL6fq5XKuPUq+oag6BgPEgZOODIMnW+8iv9lzoUbuRmJrfBCSj43KEt/klW7zKz
Dj7o49S/8TmUMv9G9WAbwOR6ptRpI49wqkE8M7eLs3zsNIZlGSyd+Gn8C+tqbv7VA/r0pmlxs8Q5
MpqvUQJY/F04Pl6L1EOfMMH08g+wcX6uoLIMGJVuYSz7rz2xNyaFpNKN38VxhOlTGbdvkWiq0HoB
Sl5zJxoQVgeP9xoDBQKF2k7g4PNL6HXWdT74vEQfhPRBWRzesAAfOt4Sq208WLzSjoYqvqlrpRbJ
OhcmWGn2rrkjH4ZEtNXOPXezekGOtvsq6yuGnU+FnA3HJiACS2vlVO08cRn3wd8KSIsmon/lSgH1
HzpNHbviZ/czmTxR9o1QZ7SZkDFAXQU+t9DS8o6KMROOIIuJsn2xiX0eihRdqldZKhKAWea6Pouy
bFllW2HZu4IC4lN6QbkShHjmWZJ4rN22OiZdNibPz+7ZLxvNh4WIXRNXfajvJCBQGjdU6ClNmklO
E/CuL4PDSSNiY9DsZ2IsdEmdzIqjdyORLqAOpWNibpcuwYNCzcwNheNimDWcOdWIvHGxxC3ias78
tAvLsiRw6P6xOIUmIGcnFxMCuopVAFMakypzZ3yI9FVj2vMw4aiT1maEq75E07GKcTqP8wpUZQmi
Y+T6ceK0zUD7zhVQu2JCIUXFEE2WoC4qPwJmL7aSotLg2F1D5wOecty0x4Save8Dabe77eH+zWsS
8vI/1zYDm9m0P0/fNL3wmn+nwRq1ILGPhAIqSUYvrTsQxT660v5DzRiqhHMZHv3xtCEpNrkScBhJ
25h1lDkGpudAhWRg2Kc/ouDREv66n2qV8rTIQxUEmLcSXbSYogqomdYtPuXz7PmMFL2ZN+ehpcx1
44orQrvqukGk6celOmkKGgpXTpbNs3MK1OeMZDmhpXOq5Sf+mjmvW+UH1zvMExUBldVZyxukGtt0
R0hg/Ti2MU16pPdKQ8dbRoCYQm4FiMb6jYFpu6PT2eHRTqmMUP2DjMpHSVUPuCULZHy3AfxTciD/
i3HfGRSKbwxljQYE+CdMqRZ/SygP5fYe0glJ8WyPl2JsemOzPCHaBrUL6NVgAxtPgHWXnp1SPiQN
97RVR0ocXqf4bvoFUkNJtvV9CWv4TL0yfTlopxdKFxebpzJaTyHdqnSPEBcSbXLaa+fGQaWBBnfS
0a2HICU1gdKS0iHAotIH9LKWjlMsHCEpAhc7ZsNMq4lObNpiitAmVLC8EclZcdtITesR0WOG4Crz
LhLwGvREt85RHqaKUF8oEIs8WNmNm1gL5feP3FumAty7C9oir4gOchKFTrhmpBGfmk+QXRJvQuuS
veR6HSCMnm86NU0UFNb+65uafL4mur/MpX1MKR+92YvWqmb98RTPTfCsDZYeThjHP74kAFonmBGR
90ZpHjIy/F1NT23Hwpc8dGLcnNRbcCrX7L4dT+wfG44J8WnJYxWQLlII4tXxiutXwNY30j+GA6RG
R+s0e1aeqUH5WnfTtpkGaqVTUmL13O29RudPVOiWM7i6KZQXmKPplAeSMUCZ2um/T4tyEDQYukVd
/pl1KoS+PXVZUWSLIi1CI0JcofVsm2ny3sBix6aMbUbBqFkl4iFxidnhh658Icsubd7vZW2bmu74
OEgZfbujUYUw3gBVcy5qnKTna7jkus0NZ8ZF09MTPwAM0sJkxnCI4tCdYxTLYdiZDSAkO69rRoP1
DatyhNaQH95WvhxEPfTeOsCPaErBHUFSgpRRmBJ2j2jCdeW26wKS46uPyLFkOlxj2uIG6TSFe3DL
MJlkDiraO5tDYRFkplRb4NvzKnShwL9ih6UZhG+wMCLnRs/Q+d1X1OzBYOedS+468ZHsMr7rTEn1
ziIYomhlhLykcMQJnIqInWy3j9CdI6mejT+IULQ9YZbAZGQYExgIgxQGsirq7wBXZqIGd1qKN8Ir
OU3QMq07aoZwyPpOqQ42V/xtMaGVGhdVL8THdXb+hSDbOkuQkHq5aysBmoDpLIoh0E4taVWuHWTD
DAe6syoxgicJOsJKQZFiItRDisc9Tto58eHFBzFubRg9t32Mr6btPAAB9AP5e6VwY+LYXWE9EW8p
BNbseqyYK8uIRG8al1kfdp2kL9dBuV0WqHygEnvjXNPXBBT/k3gJ95aHcUzm8IIRvxxN/nQeLeq7
E9UJ1m9OQgWH26UKDKICpte7fIT/bLQTVfacX6zydbD67eMAJNxJDdabEsZKjrXAR6ndnS4Opw5h
bqVlA4pdxy2p2PzxObMLuQ14LxYT54xD1PjYrolFd2KhiJ502f6526guP38BTsufla5LG/MRkAmM
MCSqUsShS6X7P2taa8EjVYV3QYG/b0KLYHUkVDOn+rss+apNcF6MN2RZrSO/Z3u+v7TZ/J/QDz0y
TNxbYhNQWb7+WuHh+QlnAGO+gF60mTHoSGu3cIuFTWEBD+8S1RFgK2zAF2Mm/9s8kISYFYAg8YAR
VIPDgqDxrtfQCmzcIlR90UaDjcpM7gEM3d/5EWSKN5vgKP/VEICo8oeXCGmMEOsICjvJWccPNT8t
rtdC2ognuRN/om8AlC9Y1OYLJF74DyX709eu8uUfIOt5cejBq29QkXuRRHeT1rivXsYMbIPOERPZ
E42HY+HQib80g4VdoykBrfAVkcqn8kILH5kBYLTlh+ZkY2XvxGnijdPCWYuj6uEAojX4OS5aB30+
J69EjdQqy+WZHGekq49ljJ9dnAopgCVXKKOsYXlH9dp/I2N6Zvh+MkImtViR1m1sdy9uxhywIJ/a
Fd4tD2c6WzXDtv7YQl7n1GzrU1lVvDamZlGYHn9FHIhnzllZClEjg9gAQhUoQRHWRX7H0T0bo6vR
yXL3oADBsu/PBKgtHWqBOOE2CtMAhkkBHK0jBYVmk1TMC6ap1A2YLNcrvF7/RMrOm4drCQz2QVM1
XJOxLQrDABCqUCD5jI8mbDVn5E6ycwxFLN0SoVTR+K2+jqLfxHGQC4/hfwthT2OMdiY/5QJhxqSN
+nK2/v4RjL5vtcVZYdQdvkoslhnrImL36WpecnwsHVEQ+aqbHHI7LIwCCi4Y8F4mqrQ1QQaBv2JD
d+jcJN3HbcPGehCaELPFgY9WwLaQf+EYAe6dp1arrxTunvTXOKzdo3ex6UnrspRdjJ3gW1HXOjAL
+oCllH0awiONj4Hp/3rlfmB28HFcTLGih+kS2J0K0c9tyNjD4UjvaSNN4OYfr73liOksHN2C42VI
7jPZC3YVAOm47HHdJeUZvq04Umxa0pcPs/OvsWV8+hYbSMsTXY1dz7C6SsiDxdZbWaDtle8hlMOi
6RY9RQQTJv0y9kUTo02k665DCoOWFpEgjxWpHIvk6B4uBiFToLGLNIFbQEyoZb8QbxGfqcERkMIZ
OX1LUIAWXwCLzvsJEvPAkh8MTbZnI39WSoJ/iJnv5B8ryc/iyJJJSwAm4Q0vEeLB3Me+x5Flx33a
MMGMy2QiAYqogETIl402/hWKJG9Gx/GwLnBBdwQl0d2QhIdNZGfv52HNxkwEmZXNxsV0K5A/By7C
ncWy6xCIGRM2QYMjGmnASUCsSkAIxncjhWb65o0bjusWihai5GQyEdtENqlXEyj7/ZPd5InhkhTR
kNISEeWzP0J9lwGU9BVofR8b5RQFZvbppv8b62YEM/Tfh41Wvvoc0cR+1XFeYiCDgADekN73nobV
P29DsvQcnXdxC0LwlhppEf5TOnGve982AqQFuuy4bOGNLu6ff8fVR5OX1TYMZJa9vYVjr8+VQzoo
UdyYkAmG7c2PQowVuI6BpUrmdQld2mQ+TVFWvJykY2jZ2yKd/duqEravshqHo19fs12te9LzlU+g
1/9XM6rW0UlU7OXp6xoXFj+0gbYX589dCAGsiVG9uPuyb1fVaYjErocfm97GDj2LWj6zbryNMw9h
0YQAbnOQiX45DYqqq4HwSonFhdDgvfFk3SZOSln915y0Wfnp446FuLjCtrbT3iQubC7hfowxCwir
wmDqNjyzO9rruZmJ4ZcVX704Ohh3ZamWA3o9LyHiQgV71+Z0B6yHIvYDZfmYC5kyoCSbqov7hxdm
gtTv782cFfinF4UfG2UR8TEkJ/WrtV8kwOTjHsNbtN1HggTZxAZ+qb49dV+rS58YEmW84FBb9EpE
N0VfkId+h26CGnQFmpRxh0u5E0j8AsezYOEfaAadQcXbeb5YV1s+S2v2EBPf/uS1RVCFOUGxl4+3
YmNqj5K0XXeONJiOV5bIMm3BAZEeoma7mNdJ4PHJN/Xgm0M5eSpgAQjz+DEYPIvaKM1wpi5iTsLt
KHkNgU6lQMizQdmgZJg129qpvAYdkqnziYeS+E8GUXg3CtQ9Lj9uc0LeM6L1TfjaXG5Cgz35HBis
Upf0gBjmflMQruwF0YJcijGdfX4ZtcmgEaCow4grGroneYTa2HIDUk3ageH0iRofv3wZ3ZYJpPO6
pUxAOhCvGCa/zf9fwU/6u1qOw765VJuR7IF06c24usWDbpx0t51URmaH0OND/pfDA3bJRHhOlwu/
L+jzZ5vo3VQ/PfxeVggbxMEaSKVClKfD5cQnhSt17WnMF2NPa+gYj226TfC/qEyJ74W9B7DNOGQ8
BCyiopk3fXzfyc6mfM7OKYxbqMoRqhxQqw2ITnJlghTyh9DrZJMDLq+q7tLjcIaiqrGf2MThnNx4
pt6kMNwGqt1EC0uiW/SWMm6OxG6bfEsVNBiR9kgSTIwhcqBbemLGMd68hLo7m6ESsnLg5HqsnDGg
K3ojEDwc9RGCjZJSXazy9D5/Zrdn5aUYFla6xkgPi9h1ACxJIhEoGgkJ0uQB0YcNPeeP14VctaMn
mVV/eB60/w2lwz6sTfz9SsdN6UrFC47+srlry/0vQq8s4pSrbfE6a0NxudJfaMfBY/10P4gLmdQ+
pq0Ve53+dFsWrzBZpRfJXgJXLckSGjkucgibighpmdEBKxN0uy8atgmKklkr/QhzurltyE1MdSmH
29hFFX1VgT/5B3RU/sdH3/ZK8qWnQW9P5d5eNkftCXymPZcpq9WtjeLzjY3l0M76f9KFmYQoXkq4
sIV9IawXddWIuOlABbxLyqbDNAddFLC+c7ht0ZcEHTYsG7ck3SR2e9gJTrEPY2yIw5NQiKgcIOKC
2rTGVvSjbKuibw1DZNPkR763lOjfCZyqiHt6kwWqBHoPbG4T4hAXSi1hwYPgMO+/7x/4hrWGcWU4
xKFfzeoEy1sesy85E3zM7NtYlH6vNc5lBq1j3CBQVXUzYykWJGe2rT/Cnisp+Bf2uEHSi8GPllH5
yb3+FZ6xHiSWWBW6akXns3TlLBpK5bMOW8K6Wn6whUg/3a3ReHUZEj7Ulna7AP1FfdJFzq0lIIsQ
+5+gUty8vUEHyDk83J8UXo31K503qtJ9zOFDP40KG1eHmaNzmWminhCejrxO09UjaHKdPJvWGYg2
u74aKkniFhcgZlrzGQqIgl3XTwCzr2lz7gk2DeO0TPOxEW2IkTV+1v33EMwbtRK+rBCyfDtFVxJs
KDz3MIEidQIHZYa+/AbbQPuW0C2A+GDQRstSXPxQ5PnWyKPBg9HrrrX+1A+zV3v6WYjxgFA2op+b
0Y14sDzcSUeyCBz5SE5eB7kwXiEOxDGdXzL40JlNvXlZ8cxmd+SI9utIWS3GUEBzlO6TGRosQrK3
Kph5oL42+oaf17pfcY9aOGH6lDwVCT5h5jtIHsMWdDa6hwww6stGnMFKP3n0MjbDKSfFg0GDAyvB
lV5lAZp6fQjvNev1T5kV+Hmsvn1pDum/3F1QVaF37cZM4hXotrWyLw4jhJ+O4M/lZx5D+Hl71BDu
H3ma+N6y4BN9hhKBifUsopadwLD6+r/wJx34x1kxnDrwk4ecRXfcf8oMLc9Z232F8q0Scy7nYsEU
TQWDoQsZJs82wtb8E3d7hTMysAhwuUyU2G1jFYUhS9yEL5T38MO730kvLBHq7HoQq9JDS9ELQJv5
eyDOSraXegvU6+cwK+F/F9l30w1LVgyfwbhA/N6H3oSuxvBH96mhXimyiHLQ7kWHAbUQfhxbNF0z
n9vcYPEv1jycug8nen8VRE6ywoEC8TkZw84dRNMmqQ6/E+9jsZt03Xfywr9GR1VSKDL0M6gsZLK5
pwjzMj5LjtRlzXzfQH00yHLaAYO95Sn9Tf5u4o4CDQCFJ6kwMIF0MEI5Srhqsiz/Ff+rbVwzwCyr
8ItPbmGbLV5ze1dZ97ggezK7+y5bqnftO74EPdtXSEC4IsVx7G78EyLHTDi8z6DGyV7M6qQuRFo6
gaybvV/EmMKefzod8BcNtTGNI63wLN2dzTgGWsl78xF+j+xDgHQpgtjTxMRsWvfMO08xpBg/k4E/
5qcib97Jpb4W75YDhjKDR73WZtv8+suF7NiXEyU0CBqrA+C6zGXJcj2VP3GF9lAF9+4pw2Uf+FO8
Iv2reWDIFbmlAhWdpjBKf0j5+AnBw1jS87zdqwpIqyicqiicQPbif/WhUgrU8JOSmxa9s4v4nFtr
tL81
`protect end_protected

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fqR67s8cBy/jbTeN196DpIBrWP6p4S7KSN05JgotCa3DCQok9PHpESJ+/YLHnMMyfVgYu3wMYulS
KP/HOuKOPw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o2f3dkiR8+1URrsaFkNAXM8HKCsrRh7Sklc6YYRJzdPn803OFcwNwVYhAiEMEOIJg1X2/T1BTFui
EQHVCIO1VCJStauI6Q8S2fTEfSbCGGuhlpfWUvhI0fluVmKgzRXGSxAPfzqyEe5IOj2rwzAzUH+w
I3b+vGSxoVxUbGLho4o=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ad3ngiL9tir1+ET0s4S3c+66wahwIoOVYNaNS7rfCSvbfk2aPsU2XB63og9D1Bg2SAX2HS1BQP3j
tM8/wIjLaDyunyJe0pY3Vy/MM/fpwDOYJVu9969hFmFD+MKjWmgclI/zBXndfn3HroxBNJ5YqbWw
T15thS0zDy/kMUmQm5Hhk2FofTiKZfDwJV8qMOs+IPoHxa32u/A5H/GAlLbYSj3iKXMDwdX1qvMx
Y/wH/Wca8f1dMVlyNgkzE7heSVl+umU4imcINE9Qacy9ksyf46mM/SkHQVg8M9UEek35LLEeFt+I
FDFYvl4xwj9zXwa6o3hy3BjN/8PdN/dXT3nHmg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
17s30izSWEvAAgQv6Vh1FDrqsfTI6ntDPxRKHcyQC5iftYo778GlTYz8H+ZoqnbRpo4Rx9iJh9p+
faDV0wcwXzKoFudL9jIBKm+gYqfFEvkVVJxOAlF/jWjG2nF/VmEXgcx03HwRaHCNUzX7tGZCK7Sm
cgQAO//GQtSMc3uUvyg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ru/nQZrQMQoFSUTnxErYixiyU4ARIhOaWewtUIoITFUVgG9z+gMss2pnsjU/kUZ9RWEI12+FXVka
+gRYtVpCxIPUEsXDftLv17WDI1tjcj5fWaceTamezhm6KUczosnGz9+NwbFG5z/2igcDAy6nQkqh
V58et0XyT53zqrn13mIfMOozEcd9PQwsZNuQCbg9wSERwoxnPdBLEg5UXNHZ0s6ahlbNehvtbbgl
yyf6RAnPelMgF4kT2YNl8xE5TPA5Ftff9vYHl3maAuj8YQ9wGLdONKEnZno1f+5yR5ljo2CbWnO+
oSovhdK1JX9QEbIkJ2QqxqDve6XKaLZUt7uHvQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NF2iKYemPHtuWn5hnoRCuPNs4c5eCM1mW9ddVILQydQ1OxFb70v0HA+tFCvBdEc/Oo23RE7HCPKv
BmrL9RcO1vKsdu91oZA6FdC/0KF7Iok4N8JN7IggHYwqedBTXbT1G79t+dcJQCYpp8IWyrFodnmv
7En+ptUiWn4gmkvJxLwkJl9miXUxtGBSTbY+MIpFl4u1hjtD6y8qRkjkITWWniMoIGON3+ShxVdH
vJ4+gC14V0VTb16Wd+kS1JZLUjkak6YQE2Y/wI+gM1SfXQv61yNCkzn4q8Fc5HhMXu8wvrAjPOoS
ZjZwz52Ph+N3YHEMsKW1FO0on8vy3THenmVVnQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4768)
`protect data_block
pa/mXep56TnCuXj5k+7cDZsyudF/BgySsJRGxM0CTQyXaSNE43YiJ69HEvLxTJm8Ea4pTJ1v9WXi
nTRcVg9K3DHOhOIzICKejreObn6KOMYE3ly/M7H+fhzllYOKD5pkQbbc9CwcFdgFf3xpYeeyEMz4
ZfzqShUQvqbeEUW+uRkz6slaIQ0IVtJMDveX3mdTJh7Xg3F17WMhx7URRVXkT7tlrfLkSDu9eN3o
+ZCIG/0/eZyjr3b8f0GIdaODojj+vIhcWigfCPa87Uy5S3/HYQpIeaD1cVEsr0wXURV6YqniErTB
x2Yz/FxZb1hpANi9M7CKVSjT6VpuBde4Fec7+wFgP/oCYh+2AgUNGVg5fM0sdhFhOQSR2bNfbr6c
PCn9CaZ/rzF6n1I3LyfCtiijML+i5tjEhSOQX3F4FtscI5PsiqCFQaEojcDWJs8NU3JpQrJuwayW
zMaq7a/1iSKj5qsPVWt/xZSkN4cODEg39klQE0U063rG4wVfrcKLF8gxWuNjw2FLsGYokMzzaFbl
XimtjmN/8jKyxl2y4zaWvxMcff/Cxw9XMvn/v4NGMs3DCrzYb7ODOT1Qbb3y5yL0X9XNM7iN4yZF
0ycB6kX4wnHmtx0D9ghdQ4pXXaIg89KXNiNaRIL2DDfbJoLnX3oXgdBVSs9GBUzaPCHXZiTDcPev
xZ11OuQSQXAI0dk79aQ0a96Z8IY4rC03j9W6wZxLJq4wVrr/6oookGD6H/5TZukc9PH8PKKjy5PE
vhzX4FIwr6TWG7kzqK+rQ0r7/AiR4vr5+L07rZ6cdqp9VcCztTi/SreYeHPCeUg8AjSdOYvU/lnI
7m+/2nWzMb0Ihx8twfJg22GRBIYFflj8JfIScwC16S572RoajOoL1IVr77TO8qdlz7rGr2zaFohr
1sXWrpp2JNy3W9y+wHkPKgjEpmVSy1+dFhKdl4ZZkiJqHcmM9EgbtC28iRfl8PQxaLKrbcvsRjDm
ZmYxHdqlesZro3kuS5Z30Llj+N78aWMYFpm12Wd30wA/WiTY0g1nzO0NJmOMaHW6uU1Bp8e+oTKu
gmAjeWADyVeBnhsdfgoGUkZlN6qw73EOprw63IKrKoNu6+W5jD4CaX8nEOghL7NxLPO1yohOBnn4
zvD9ZKm8XEl8N6BoqupG/FABKx9evCsqMfbr6xbVDNU3O1KMJXvToPedonAy5GfxLJKXk8mQxXCl
jXcmmlhe3lVEiuOukxF6eYYYVVcT5/oYLcchlabmKyFZ4x7uKmA7zyev/CnQPhWvvN48Z+s4Rrlt
mI1Dgk+YrJ1zmQAkMFKOWVQqBsyvydZT2n562MGT8VDN0QgrlDfs9XPJuK/biW6RE59e0irs3kB7
w4IOqfxMK5qlVLkhBmd00ZJDuNOK/GdhSQNxJ8A8RtF9cBfsqMbHCJCYwCRJMUUBk7s1QfeSVuaj
StEW2+jNvsi7oIR0NWjJgUWeqkbO5QQOma0nrjgwoXwlCGQ4ouVDQj3dU531RH/FaNIgZcDKRFtA
Nbqzp3ofNc66eiIEY/CP0Xh/a5CCNbu4BSwFrhnTsA3knTbK/o2bvMyFsqgCZeuf8TJai/H/Ol50
9meqz3gTueLV0F75aq/CbGaTEH+QhM12UQPnUPb7DQWx/5k7eSSuYZwnIROQUj7ZBX+GkeEz7oOj
4EctmgulZt8P5zt48i9H9NW7OXsKLsKgFMa6lAAgrGKBlFwm3+jSQb1kor3canz0JFRQ3tE8FCRu
aZc5Q4K3L5nK/bj79/n9zdfehcpX6b0UYqolsor2LkQvHRhzX+vu79BRcUN4JKPqp9wBYf93YSAQ
JnbcC0JzPFh/l+oI6YhWcXOgNoQWoncHt/3qaMfc50EiGiK3vuuht3HX3923RfpTC+0DYjCP6LVO
9GnRZAQiwSEZ1jrm04kj6n1c5aIKvzzz9s6CYPv53tf2YK7ZOFg5PO6ucZjj6NRkmgF1IrTa1pBT
QTdYgBUqRydD2uTnlpW5LSvxZy/Z133+kTPEz9N/rY4ZSYESk3c9OxrHbHGUyAvBeK+hcVM2I37f
W4MCo2d9JAu3vlleFdae8BD8yaCmDqf+dGE0P5U2aY61hh1SLmg0OyRv9CiLdEphjPYZjnJHKyRK
rmLA/c22lsSAcj1OIwQXd93qxzngiB8uckZWL8EZ1hpBO4xgPLVsEePF8KlVFkciLnX8aQkkTc0P
DDrh3OT/vQMgA8zK1EHrAjNzevTwoWJJNOhv9D+Oe0AssNlByBNxE9kDZ214o0V9WQIX4vYCt5Vp
eEvbIKmQh/rl8DTswTHE5L7FbXPZqONAE/ma3iCG7nlVLBUBg7WtjgJ8B1o6KTDMSZI/iq2nF1w/
D5e4w9FLYQ6BOLtQ1TXzej4DKqqwEAhzDtpKFpDTMuthykjDpMzOwU2esud7XxiebHbL6xFBix8r
w0bT+SQyuvoXGWzsDOxnzsOFuKXruPqfmJAiJvlFeV8GEQzHn62xw8QRwkaPVgdd40bmBv4D78eb
/vadY4msjk2e2WEgXgPxz0W3Iw+uTbf7aFBaWCmmq/wgbve8XF7+qGKSJTKbxFfwI+xtqm3ypVUJ
U4X03E0YgMqQ5GphPEyHrfdKf4VFfkJyII0ebPmIHdH5Kq1/BACS12NgOco5x4DAH36bhTHmykt2
c/HVYw+n3+TjH2bKjd1A9nfeqnDVhcmGyDnx7xqafX357Xb4AIZkBU3+XJ8Td1BAOB0jckpFNgNF
ohH8EHWHneLiEuCXZ2odiMFL4cnmRSMypNX+2dF4EX3WqYunGcXpDzrC+6QtH81qg7O7Xc+uxFqc
Z/yJ5TPc6f1iYTMnd2Xm86oMUmr90cLr9Nw1uHp2mpFu/W2Pv6vBPKZYtXUSbe9cDllucnN/ed9s
0FZwe/Az88jvXyAH476A7+23DTo0LtPdmEfJmfwl+OBgnKMIIORUsyGRKBzwF85dnkg8Pd0H5g02
IZYgZCxpz6HM2J7+zXS7ZiGFAvaGDasqytVOku6uCLwb9vE1MKS+aGi5zE0b5QmofQe4+d+Po71H
h9GW0kVOtQJPWOYmL01IeEOIm7dABmz+SipX1XIsfekcQ6V2/pH6tD4MTg+093L1Jn5fWnlit1Ku
JlR3EQDoJTbooYhcJEISeUGqeSqvDquUN27qXBMUBvCOunu/BBaw14ueIXBXNz26s5kS3T80k71K
uApu+Gk4j5tkeiQpKy8htEuzfBWn1P5vvTSDk+QpofxCOoRg8lQ7HodIQCirUnjCmHFWF+mbhbeK
dngqisSVaLVvmjf0A8DTH+ojy/62u1jTIvZ+agk/N91YVAJKhnATE/ctTtvhyYO1D7jW+PQ55wfK
5QRBducZ4JkRCGoqQEiqdQC8yTZEza547n9z/u3VX71bFO+1lfR67hj+J1h1MMsox9hOkFiEU/h/
b50hOhkdZ0rL+asRC8xosm2DUtjlnN5UFQIvqjg+5YWxuP+8g5Ddrxp30JCPb87WXjF89bAGqsz6
GCKy1V0xE3VjP97u1+OATkjrzyjA4Ge+1LOyzfLMiieT6ARY0w6zi2TNk3TmTQAFYrVWTnHfWdsf
W40+XJrK4465jWBgsF72lM0I53A5tuEPvIHgo4aSckt5gmXQOZPqGlMfpzDMBC/lh0wFQTTCU0wc
661SsKDCztWyuX4lkrRZiqQ2OTgBjGmXXjo4PErPUpyBhDtvH4548d+iN3SdRG2jgX3qHDVE4Vwr
Kk8eATrnHrQADZJTWbqaBzKvG0T383KsInnpOJtZNAc3gWbrZyRU1m7Lt8BJq+gzwnm+80PB1Vb2
WntkfBFyqQLhUiqqEZ5CLPizRTJOMMCZd8tVLp4aEwWvKd3J/HL/GV00zzkUQYxDYljkwkMHueY2
HqH78QdBhozJOH1cga/fwjLd+CArG+Nr+K6bikIn3gDelYFhvWWge2qaXN+MeuGC7xJTaXSSiwVB
kGBdYbL0XsclPd07NPOTyTQI5V7toMKZp241oEeIrRdo+LMzyilZIZ6Kc7eOGG4K6A6OJn6QFAdr
p7UOwXQkaZZl016IgpcRA7cyBwlbwmJd7DIVZY5pONkWZl5+NpQf829K9rBRzJ9b31fnj2TcZOR1
3wBxK8z9XzePmiNTMRmIT32t9LYzTmT5YglLIGOgErZBnoae+I/Q+SKKBxRc3Xe/AEl3x14IBHhJ
urXt4mpEysh2rwWrrTuVCkuHH3J6iUYDDYNyDsH4nClGN5axVjhB38WqbsjvnXTz9QbEny1O0s1L
R6EGlrIkF40mVj2sN+aMdGnwnIXLY4aZ7lqMnA6EsiL8icFH8vdLJzXLwsZWezw4VCt2X1Jidi6/
8Ssv8ycCCgC6bDE0Wz5NUzisDwHi1jSNgHwGTPlZgYZt28U4dL/lepjByKe944CZ7/wi0i/rk/An
tafpU5grwzSXpBOShrgWLN1xf8qbCPq2ul8IrHdo/mfHslocI06yJAGYIsqXaNfHVumHEEQjV15g
8kmNfGhzbMrDhWzqvXityr54f4JOQH4o4Bbpr25wvM3kbvy+WaiCOuUVr4YE5DqQIRtt35XIJO+2
XUeAJk27OECNIXP2fVYLuUj1m+bkWP0pSZD/EXfueIMvvs5m5l/gXR8x1E9Rqb15Y/d0plGEdNqs
gZDvDOAFEwlgxprnlcV7VfRtHib1rLCnlp3SRRxYOhcPz2MRdRfgOGnz2Y2KpK429TfwKDVAFFkX
He0UbzlbJOK8YskgYy6Qtm2WCM8ukJev4cqs4jD7nYy+C/1shtCXw5Z+XYVjBHvcZnMHnon5cHSp
UcxClKzkABD6Ah5nNPsTXNubbE5WVbO3erESEa9okxDLyJSkR9DyMmGcDU7sqAS2I/CZyGNhHdWH
poeWFPMMi8yP219B9bBfKM8wXfI17bTD0VS8SBN0LcPu8gBOboZtZc3NVYNxjiga3Uluckfd+DrV
Simr/rAAnlMmSG7c66GsVMj81N8MGJdMdGjANR5S/yLW9Lr66ZCTN3y2E/7AyIztHqmPLwt3K3oM
gZxtCcqgWocIknBPmxf3kF7KLbnceDsxKGq2HRmvvQjgH4SUUkk7Sm2FOIRtLVAxhsjxeJW2HRbF
g0SYJSaZg90rd7nYBC1iOqg0PrRh1gkb0rYTrMvb4Ee9dH5QEGSGrS6gjQ8gH509apxilMJLgPaF
6u7VLxkZWxcsFouw/E9bqguBtcjhQaelukA9L21ARvaGQ2UXC+e1eyjalt0XLgJK1dnV9Rt5BzXo
qgpJ4axLqvxT3cwQrXhPfu4EBS81triMNbpg4NFYeruwt34w896WxI/+ETl+uFYS7vUx4H4i7gd0
TH1ciOPNBWdXkicdx9poB1zt7oD+vyjPcrl77/NrF9I2wRU+m8FfZKUP9QXQCCsYr2tvP6dpbnY8
eIxTnXcxelO/IUKH3gBn6zcHpTTWw/7i0DOJoqdYayrACtpt1YjxzzQx//Clv6ujQpOo/JEIXpWU
GgErSNMR/ZWZrzZGL95lg/MYdAAkaUKejlseCQnDVtJmAJOhofZKjpsrnQeAMcrDJK8QNsn5ZVZv
Awy6gEjEahxKc0kkvQMhIBsjhnSDiIVeIyr4MIEPCn11pgugX/oSU0JUDaykcU/t4hj0v31f7Hnq
FlMsWadW9/zTWIBbWDBMFZU2yqsrpn0aCStn654yl8y2nQPJUEgdbx+T6u+aD6INOijCAztgNL9b
dtg5B0r4JQHZtP0waVkhbUnYJeDRU5JtryhkX6WgNled5WdJO+hupGJDpnEJXoK5MY6fI5JZDqiM
zd01L44Tjl1TSHBINv8xU6hyPHpzipnOjVoYBxrHnUp/8S7krYcl4d2roL1wHhZuBXl3wT1pZ+oK
ksFtJvoCIe83z1lj6N20fRuJrIiH8+PddkiQMfi6iYm6gHBMJSUkESULQQ1hyqnkrDVLjXmtlGuX
xkDbZZJyMGdlkwlEhMqvg8YUSHO0tQ2JaSmIgifA5aSsC4Tye0A2g+WL9dtTmlaSZ7sqyj6G+mLf
JhdgNyvNmF7t0/QD57fAmyVSQvNLuDQ0haqq1Bli4aD35ST/UJ3KdjYRBBD4YNrRXlRyNv6rx4tz
z1WYaQOLrsy2hl8In3HcdFY3EdzXkcAaaI4ocwNRv/+QJ+GJJdoid7YVtgI1KBPqzobkWu10dzuo
SKMoxUMjGLqIcZ/rqnp4+qKiaXwCCNv+/v3rMCHXIjrarGkwsMDL9DQRPePI2UJgwtsfPbLoskHT
Eaik0gEU3R4Jvylzi0jAg1+2UIHAsAIsEgbMlsIF5SpYUm66Btx0wQA8r8UQgvlRAEMv/dPaoo8d
DuPRdjMM5oe0CNlEq5BT1a+RDgyiOJm/jeqQpq662gozL5bBrw==
`protect end_protected
